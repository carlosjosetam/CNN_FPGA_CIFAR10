mgc_hls.BLOCK_1R1W_RBW(rtl) :16: :11: :1728:
mgc_hls.mgc_io_sync_v2(beh) :0:
