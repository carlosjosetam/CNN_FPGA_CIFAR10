
//------> /softl3/catapultc10_1b/Mgc_home/pkgs/siflibs/ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> /softl3/catapultc10_1b/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /softl3/catapultc10_1b/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.v 
// Block 1R1W Read Before Write RAM with common clock
module BLOCK_1R1W_RBW
#(
parameter data_width = 8,
parameter addr_width = 7,
parameter depth = 128
)(
	radr, wadr, d, we, re, clk, q
);

	input [addr_width-1:0] radr;
	input [addr_width-1:0] wadr;
	input [data_width-1:0] d;
	input we;
	input re;
	input clk;
	output[data_width-1:0] q;

	reg [data_width-1:0] q;

	(* ram_style = "block" *)
	reg [data_width-1:0] mem [depth-1:0];// synthesis syn_ramstyle="block_ram"
	//pragma attribute mem block_ram true
		
	always @(posedge clk) begin
		if (we) begin
			mem[wadr] <= d; // Write port
		end
		if (re) begin
			q <= mem[radr] ; // read port
		end
	end

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.1b/747384 Production Release
//  HLS Date:       Wed Nov  1 10:26:06 PDT 2017
// 
//  Generated by:   xph3sei710@ocaepc56
//  Generated date: Fri Jan 25 10:40:08 2019
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_11_1728_12_gen
// ------------------------------------------------------------------


module CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_11_1728_12_gen (
  we, d, wadr, re, q, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d
);
  output we;
  output [15:0] d;
  output [10:0] wadr;
  output re;
  input [15:0] q;
  output [10:0] radr;
  input [10:0] radr_d;
  input [10:0] wadr_d;
  input [15:0] d_d;
  input we_d;
  input re_d;
  output [15:0] q_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (we_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign re = (re_d);
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_11_1728_11_gen
// ------------------------------------------------------------------


module CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_11_1728_11_gen (
  we, d, wadr, re, q, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d
);
  output we;
  output [15:0] d;
  output [10:0] wadr;
  output re;
  input [15:0] q;
  output [10:0] radr;
  input [10:0] radr_d;
  input [10:0] wadr_d;
  input [15:0] d_d;
  input we_d;
  input re_d;
  output [15:0] q_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (we_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign re = (re_d);
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_4_10_9_gen
// ------------------------------------------------------------------


module CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_4_10_9_gen (
  re, q, radr, radr_d, re_d, q_d
);
  output re;
  input [15:0] q;
  output [3:0] radr;
  input [3:0] radr_d;
  input re_d;
  output [15:0] q_d;



  // Interconnect Declarations for Component Instantiations 
  assign re = (re_d);
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1800_8_gen
// ------------------------------------------------------------------


module CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1800_8_gen (
  re, q, radr, radr_d, re_d, q_d
);
  output re;
  input [15:0] q;
  output [10:0] radr;
  input [10:0] radr_d;
  input re_d;
  output [15:0] q_d;



  // Interconnect Declarations for Component Instantiations 
  assign re = (re_d);
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_5_20_7_gen
// ------------------------------------------------------------------


module CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_5_20_7_gen (
  re, q, radr, radr_d, re_d, q_d
);
  output re;
  input [15:0] q;
  output [4:0] radr;
  input [4:0] radr_d;
  input re_d;
  output [15:0] q_d;



  // Interconnect Declarations for Component Instantiations 
  assign re = (re_d);
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_13_5760_6_gen
// ------------------------------------------------------------------


module CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_13_5760_6_gen (
  re, q, radr, radr_d, re_d, q_d
);
  output re;
  input [15:0] q;
  output [12:0] radr;
  input [12:0] radr_d;
  input re_d;
  output [15:0] q_d;



  // Interconnect Declarations for Component Instantiations 
  assign re = (re_d);
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_5_32_5_gen
// ------------------------------------------------------------------


module CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_5_32_5_gen (
  re, q, radr, radr_d, re_d, q_d
);
  output re;
  input [15:0] q;
  output [4:0] radr;
  input [4:0] radr_d;
  input re_d;
  output [15:0] q_d;



  // Interconnect Declarations for Component Instantiations 
  assign re = (re_d);
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_15_18432_4_gen
// ------------------------------------------------------------------


module CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_15_18432_4_gen (
  re, q, radr, radr_d, re_d, q_d
);
  output re;
  input [15:0] q;
  output [14:0] radr;
  input [14:0] radr_d;
  input re_d;
  output [15:0] q_d;



  // Interconnect Declarations for Component Instantiations 
  assign re = (re_d);
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_6_64_3_gen
// ------------------------------------------------------------------


module CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_6_64_3_gen (
  re, q, radr, radr_d, re_d, q_d
);
  output re;
  input [15:0] q;
  output [5:0] radr;
  input [5:0] radr_d;
  input re_d;
  output [15:0] q_d;



  // Interconnect Declarations for Component Instantiations 
  assign re = (re_d);
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1728_2_gen
// ------------------------------------------------------------------


module CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1728_2_gen (
  re, q, radr, radr_d, re_d, q_d
);
  output re;
  input [15:0] q;
  output [10:0] radr;
  input [10:0] radr_d;
  input re_d;
  output [15:0] q_d;



  // Interconnect Declarations for Component Instantiations 
  assign re = (re_d);
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1728_1_gen
// ------------------------------------------------------------------


module CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1728_1_gen (
  re, q, radr, radr_d, re_d, q_d
);
  output re;
  input [15:0] q;
  output [10:0] radr;
  input [10:0] radr_d;
  input re_d;
  output [15:0] q_d;



  // Interconnect Declarations for Component Instantiations 
  assign re = (re_d);
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    CNN_main_simple_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module CNN_main_simple_core_core_fsm (
  clk, rst, fsm_output, INIT_I_C_1_tr0, INIT_J_C_0_tr0, INIT_L_C_0_tr0, FOR_B_C_1_tr0,
      FOR_A_C_0_tr0, FOR_I_C_2_tr0, FOR_J_C_0_tr0, FOR_K_C_0_tr0, BIAS_I_C_2_tr0,
      BIAS_J_C_0_tr0, FOR_L_C_0_tr0, FOR_A_1_C_1_tr0, FOR_B_1_C_1_tr0, FOR_I_1_C_1_tr0,
      FOR_J_1_C_1_tr0, FOR_K_1_C_0_tr0, INIT_I_1_C_1_tr0, INIT_J_1_C_0_tr0, INIT_L_1_C_0_tr0,
      FOR_B_2_C_1_tr0, FOR_A_2_C_0_tr0, FOR_I_2_C_2_tr0, FOR_J_2_C_0_tr0, FOR_K_2_C_0_tr0,
      BIAS_I_1_C_2_tr0, BIAS_J_1_C_0_tr0, FOR_L_1_C_0_tr0, FOR_A_3_C_1_tr0, FOR_B_3_C_1_tr0,
      FOR_I_3_C_1_tr0, FOR_J_3_C_1_tr0, FOR_K_3_C_0_tr0, INIT_I_2_C_1_tr0, INIT_J_2_C_0_tr0,
      INIT_L_2_C_0_tr0, FOR_B_4_C_1_tr0, FOR_A_4_C_0_tr0, FOR_I_4_C_2_tr0, FOR_J_4_C_0_tr0,
      FOR_K_4_C_0_tr0, BIAS_I_2_C_2_tr0, BIAS_J_2_C_0_tr0, FOR_L_2_C_0_tr0, FOR_A_5_C_1_tr0,
      FOR_B_5_C_1_tr0, FOR_I_5_C_1_tr0, FOR_J_5_C_1_tr0, FOR_K_5_C_0_tr0, FOR_K_6_C_2_tr0,
      FOR_J_6_C_0_tr0, FOR_I_6_C_0_tr0, FOR_K_7_C_1_tr0, FOR_J_7_C_1_tr0, for_C_0_tr0
);
  input clk;
  input rst;
  output [91:0] fsm_output;
  reg [91:0] fsm_output;
  input INIT_I_C_1_tr0;
  input INIT_J_C_0_tr0;
  input INIT_L_C_0_tr0;
  input FOR_B_C_1_tr0;
  input FOR_A_C_0_tr0;
  input FOR_I_C_2_tr0;
  input FOR_J_C_0_tr0;
  input FOR_K_C_0_tr0;
  input BIAS_I_C_2_tr0;
  input BIAS_J_C_0_tr0;
  input FOR_L_C_0_tr0;
  input FOR_A_1_C_1_tr0;
  input FOR_B_1_C_1_tr0;
  input FOR_I_1_C_1_tr0;
  input FOR_J_1_C_1_tr0;
  input FOR_K_1_C_0_tr0;
  input INIT_I_1_C_1_tr0;
  input INIT_J_1_C_0_tr0;
  input INIT_L_1_C_0_tr0;
  input FOR_B_2_C_1_tr0;
  input FOR_A_2_C_0_tr0;
  input FOR_I_2_C_2_tr0;
  input FOR_J_2_C_0_tr0;
  input FOR_K_2_C_0_tr0;
  input BIAS_I_1_C_2_tr0;
  input BIAS_J_1_C_0_tr0;
  input FOR_L_1_C_0_tr0;
  input FOR_A_3_C_1_tr0;
  input FOR_B_3_C_1_tr0;
  input FOR_I_3_C_1_tr0;
  input FOR_J_3_C_1_tr0;
  input FOR_K_3_C_0_tr0;
  input INIT_I_2_C_1_tr0;
  input INIT_J_2_C_0_tr0;
  input INIT_L_2_C_0_tr0;
  input FOR_B_4_C_1_tr0;
  input FOR_A_4_C_0_tr0;
  input FOR_I_4_C_2_tr0;
  input FOR_J_4_C_0_tr0;
  input FOR_K_4_C_0_tr0;
  input BIAS_I_2_C_2_tr0;
  input BIAS_J_2_C_0_tr0;
  input FOR_L_2_C_0_tr0;
  input FOR_A_5_C_1_tr0;
  input FOR_B_5_C_1_tr0;
  input FOR_I_5_C_1_tr0;
  input FOR_J_5_C_1_tr0;
  input FOR_K_5_C_0_tr0;
  input FOR_K_6_C_2_tr0;
  input FOR_J_6_C_0_tr0;
  input FOR_I_6_C_0_tr0;
  input FOR_K_7_C_1_tr0;
  input FOR_J_7_C_1_tr0;
  input for_C_0_tr0;


  // FSM State Type Declaration for CNN_main_simple_core_core_fsm_1
  parameter
    core_rlp_C_0 = 7'd0,
    core_rlp_C_1 = 7'd1,
    main_C_0 = 7'd2,
    INIT_I_C_0 = 7'd3,
    INIT_I_C_1 = 7'd4,
    INIT_J_C_0 = 7'd5,
    INIT_L_C_0 = 7'd6,
    FOR_B_C_0 = 7'd7,
    FOR_B_C_1 = 7'd8,
    FOR_A_C_0 = 7'd9,
    FOR_I_C_0 = 7'd10,
    FOR_I_C_1 = 7'd11,
    FOR_I_C_2 = 7'd12,
    FOR_J_C_0 = 7'd13,
    FOR_K_C_0 = 7'd14,
    BIAS_I_C_0 = 7'd15,
    BIAS_I_C_1 = 7'd16,
    BIAS_I_C_2 = 7'd17,
    BIAS_J_C_0 = 7'd18,
    FOR_L_C_0 = 7'd19,
    FOR_J_1_C_0 = 7'd20,
    FOR_I_1_C_0 = 7'd21,
    FOR_A_1_C_0 = 7'd22,
    FOR_A_1_C_1 = 7'd23,
    FOR_B_1_C_0 = 7'd24,
    FOR_B_1_C_1 = 7'd25,
    FOR_I_1_C_1 = 7'd26,
    FOR_J_1_C_1 = 7'd27,
    FOR_K_1_C_0 = 7'd28,
    INIT_I_1_C_0 = 7'd29,
    INIT_I_1_C_1 = 7'd30,
    INIT_J_1_C_0 = 7'd31,
    INIT_L_1_C_0 = 7'd32,
    FOR_B_2_C_0 = 7'd33,
    FOR_B_2_C_1 = 7'd34,
    FOR_A_2_C_0 = 7'd35,
    FOR_I_2_C_0 = 7'd36,
    FOR_I_2_C_1 = 7'd37,
    FOR_I_2_C_2 = 7'd38,
    FOR_J_2_C_0 = 7'd39,
    FOR_K_2_C_0 = 7'd40,
    BIAS_I_1_C_0 = 7'd41,
    BIAS_I_1_C_1 = 7'd42,
    BIAS_I_1_C_2 = 7'd43,
    BIAS_J_1_C_0 = 7'd44,
    FOR_L_1_C_0 = 7'd45,
    FOR_J_3_C_0 = 7'd46,
    FOR_I_3_C_0 = 7'd47,
    FOR_A_3_C_0 = 7'd48,
    FOR_A_3_C_1 = 7'd49,
    FOR_B_3_C_0 = 7'd50,
    FOR_B_3_C_1 = 7'd51,
    FOR_I_3_C_1 = 7'd52,
    FOR_J_3_C_1 = 7'd53,
    FOR_K_3_C_0 = 7'd54,
    INIT_I_2_C_0 = 7'd55,
    INIT_I_2_C_1 = 7'd56,
    INIT_J_2_C_0 = 7'd57,
    INIT_L_2_C_0 = 7'd58,
    FOR_B_4_C_0 = 7'd59,
    FOR_B_4_C_1 = 7'd60,
    FOR_A_4_C_0 = 7'd61,
    FOR_I_4_C_0 = 7'd62,
    FOR_I_4_C_1 = 7'd63,
    FOR_I_4_C_2 = 7'd64,
    FOR_J_4_C_0 = 7'd65,
    FOR_K_4_C_0 = 7'd66,
    BIAS_I_2_C_0 = 7'd67,
    BIAS_I_2_C_1 = 7'd68,
    BIAS_I_2_C_2 = 7'd69,
    BIAS_J_2_C_0 = 7'd70,
    FOR_L_2_C_0 = 7'd71,
    FOR_J_5_C_0 = 7'd72,
    FOR_I_5_C_0 = 7'd73,
    FOR_A_5_C_0 = 7'd74,
    FOR_A_5_C_1 = 7'd75,
    FOR_B_5_C_0 = 7'd76,
    FOR_B_5_C_1 = 7'd77,
    FOR_I_5_C_1 = 7'd78,
    FOR_J_5_C_1 = 7'd79,
    FOR_K_5_C_0 = 7'd80,
    FOR_K_6_C_0 = 7'd81,
    FOR_K_6_C_1 = 7'd82,
    FOR_K_6_C_2 = 7'd83,
    FOR_J_6_C_0 = 7'd84,
    FOR_I_6_C_0 = 7'd85,
    FOR_J_7_C_0 = 7'd86,
    FOR_K_7_C_0 = 7'd87,
    FOR_K_7_C_1 = 7'd88,
    FOR_J_7_C_1 = 7'd89,
    for_C_0 = 7'd90,
    main_C_1 = 7'd91;

  reg [6:0] state_var;
  reg [6:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : CNN_main_simple_core_core_fsm_1
    case (state_var)
      core_rlp_C_1 : begin
        fsm_output = 92'b10;
        state_var_NS = main_C_0;
      end
      main_C_0 : begin
        fsm_output = 92'b100;
        state_var_NS = INIT_I_C_0;
      end
      INIT_I_C_0 : begin
        fsm_output = 92'b1000;
        state_var_NS = INIT_I_C_1;
      end
      INIT_I_C_1 : begin
        fsm_output = 92'b10000;
        if ( INIT_I_C_1_tr0 ) begin
          state_var_NS = INIT_J_C_0;
        end
        else begin
          state_var_NS = INIT_I_C_0;
        end
      end
      INIT_J_C_0 : begin
        fsm_output = 92'b100000;
        if ( INIT_J_C_0_tr0 ) begin
          state_var_NS = INIT_L_C_0;
        end
        else begin
          state_var_NS = INIT_I_C_0;
        end
      end
      INIT_L_C_0 : begin
        fsm_output = 92'b1000000;
        if ( INIT_L_C_0_tr0 ) begin
          state_var_NS = FOR_B_C_0;
        end
        else begin
          state_var_NS = INIT_I_C_0;
        end
      end
      FOR_B_C_0 : begin
        fsm_output = 92'b10000000;
        state_var_NS = FOR_B_C_1;
      end
      FOR_B_C_1 : begin
        fsm_output = 92'b100000000;
        if ( FOR_B_C_1_tr0 ) begin
          state_var_NS = FOR_A_C_0;
        end
        else begin
          state_var_NS = FOR_B_C_0;
        end
      end
      FOR_A_C_0 : begin
        fsm_output = 92'b1000000000;
        if ( FOR_A_C_0_tr0 ) begin
          state_var_NS = FOR_I_C_0;
        end
        else begin
          state_var_NS = FOR_B_C_0;
        end
      end
      FOR_I_C_0 : begin
        fsm_output = 92'b10000000000;
        state_var_NS = FOR_I_C_1;
      end
      FOR_I_C_1 : begin
        fsm_output = 92'b100000000000;
        state_var_NS = FOR_I_C_2;
      end
      FOR_I_C_2 : begin
        fsm_output = 92'b1000000000000;
        if ( FOR_I_C_2_tr0 ) begin
          state_var_NS = FOR_J_C_0;
        end
        else begin
          state_var_NS = FOR_B_C_0;
        end
      end
      FOR_J_C_0 : begin
        fsm_output = 92'b10000000000000;
        if ( FOR_J_C_0_tr0 ) begin
          state_var_NS = FOR_K_C_0;
        end
        else begin
          state_var_NS = FOR_B_C_0;
        end
      end
      FOR_K_C_0 : begin
        fsm_output = 92'b100000000000000;
        if ( FOR_K_C_0_tr0 ) begin
          state_var_NS = BIAS_I_C_0;
        end
        else begin
          state_var_NS = FOR_B_C_0;
        end
      end
      BIAS_I_C_0 : begin
        fsm_output = 92'b1000000000000000;
        state_var_NS = BIAS_I_C_1;
      end
      BIAS_I_C_1 : begin
        fsm_output = 92'b10000000000000000;
        state_var_NS = BIAS_I_C_2;
      end
      BIAS_I_C_2 : begin
        fsm_output = 92'b100000000000000000;
        if ( BIAS_I_C_2_tr0 ) begin
          state_var_NS = BIAS_J_C_0;
        end
        else begin
          state_var_NS = BIAS_I_C_0;
        end
      end
      BIAS_J_C_0 : begin
        fsm_output = 92'b1000000000000000000;
        if ( BIAS_J_C_0_tr0 ) begin
          state_var_NS = FOR_L_C_0;
        end
        else begin
          state_var_NS = BIAS_I_C_0;
        end
      end
      FOR_L_C_0 : begin
        fsm_output = 92'b10000000000000000000;
        if ( FOR_L_C_0_tr0 ) begin
          state_var_NS = FOR_J_1_C_0;
        end
        else begin
          state_var_NS = FOR_B_C_0;
        end
      end
      FOR_J_1_C_0 : begin
        fsm_output = 92'b100000000000000000000;
        state_var_NS = FOR_I_1_C_0;
      end
      FOR_I_1_C_0 : begin
        fsm_output = 92'b1000000000000000000000;
        state_var_NS = FOR_A_1_C_0;
      end
      FOR_A_1_C_0 : begin
        fsm_output = 92'b10000000000000000000000;
        state_var_NS = FOR_A_1_C_1;
      end
      FOR_A_1_C_1 : begin
        fsm_output = 92'b100000000000000000000000;
        if ( FOR_A_1_C_1_tr0 ) begin
          state_var_NS = FOR_B_1_C_0;
        end
        else begin
          state_var_NS = FOR_A_1_C_0;
        end
      end
      FOR_B_1_C_0 : begin
        fsm_output = 92'b1000000000000000000000000;
        state_var_NS = FOR_B_1_C_1;
      end
      FOR_B_1_C_1 : begin
        fsm_output = 92'b10000000000000000000000000;
        if ( FOR_B_1_C_1_tr0 ) begin
          state_var_NS = FOR_I_1_C_1;
        end
        else begin
          state_var_NS = FOR_A_1_C_0;
        end
      end
      FOR_I_1_C_1 : begin
        fsm_output = 92'b100000000000000000000000000;
        if ( FOR_I_1_C_1_tr0 ) begin
          state_var_NS = FOR_J_1_C_1;
        end
        else begin
          state_var_NS = FOR_I_1_C_0;
        end
      end
      FOR_J_1_C_1 : begin
        fsm_output = 92'b1000000000000000000000000000;
        if ( FOR_J_1_C_1_tr0 ) begin
          state_var_NS = FOR_K_1_C_0;
        end
        else begin
          state_var_NS = FOR_J_1_C_0;
        end
      end
      FOR_K_1_C_0 : begin
        fsm_output = 92'b10000000000000000000000000000;
        if ( FOR_K_1_C_0_tr0 ) begin
          state_var_NS = INIT_I_1_C_0;
        end
        else begin
          state_var_NS = FOR_J_1_C_0;
        end
      end
      INIT_I_1_C_0 : begin
        fsm_output = 92'b100000000000000000000000000000;
        state_var_NS = INIT_I_1_C_1;
      end
      INIT_I_1_C_1 : begin
        fsm_output = 92'b1000000000000000000000000000000;
        if ( INIT_I_1_C_1_tr0 ) begin
          state_var_NS = INIT_J_1_C_0;
        end
        else begin
          state_var_NS = INIT_I_1_C_0;
        end
      end
      INIT_J_1_C_0 : begin
        fsm_output = 92'b10000000000000000000000000000000;
        if ( INIT_J_1_C_0_tr0 ) begin
          state_var_NS = INIT_L_1_C_0;
        end
        else begin
          state_var_NS = INIT_I_1_C_0;
        end
      end
      INIT_L_1_C_0 : begin
        fsm_output = 92'b100000000000000000000000000000000;
        if ( INIT_L_1_C_0_tr0 ) begin
          state_var_NS = FOR_B_2_C_0;
        end
        else begin
          state_var_NS = INIT_I_1_C_0;
        end
      end
      FOR_B_2_C_0 : begin
        fsm_output = 92'b1000000000000000000000000000000000;
        state_var_NS = FOR_B_2_C_1;
      end
      FOR_B_2_C_1 : begin
        fsm_output = 92'b10000000000000000000000000000000000;
        if ( FOR_B_2_C_1_tr0 ) begin
          state_var_NS = FOR_A_2_C_0;
        end
        else begin
          state_var_NS = FOR_B_2_C_0;
        end
      end
      FOR_A_2_C_0 : begin
        fsm_output = 92'b100000000000000000000000000000000000;
        if ( FOR_A_2_C_0_tr0 ) begin
          state_var_NS = FOR_I_2_C_0;
        end
        else begin
          state_var_NS = FOR_B_2_C_0;
        end
      end
      FOR_I_2_C_0 : begin
        fsm_output = 92'b1000000000000000000000000000000000000;
        state_var_NS = FOR_I_2_C_1;
      end
      FOR_I_2_C_1 : begin
        fsm_output = 92'b10000000000000000000000000000000000000;
        state_var_NS = FOR_I_2_C_2;
      end
      FOR_I_2_C_2 : begin
        fsm_output = 92'b100000000000000000000000000000000000000;
        if ( FOR_I_2_C_2_tr0 ) begin
          state_var_NS = FOR_J_2_C_0;
        end
        else begin
          state_var_NS = FOR_B_2_C_0;
        end
      end
      FOR_J_2_C_0 : begin
        fsm_output = 92'b1000000000000000000000000000000000000000;
        if ( FOR_J_2_C_0_tr0 ) begin
          state_var_NS = FOR_K_2_C_0;
        end
        else begin
          state_var_NS = FOR_B_2_C_0;
        end
      end
      FOR_K_2_C_0 : begin
        fsm_output = 92'b10000000000000000000000000000000000000000;
        if ( FOR_K_2_C_0_tr0 ) begin
          state_var_NS = BIAS_I_1_C_0;
        end
        else begin
          state_var_NS = FOR_B_2_C_0;
        end
      end
      BIAS_I_1_C_0 : begin
        fsm_output = 92'b100000000000000000000000000000000000000000;
        state_var_NS = BIAS_I_1_C_1;
      end
      BIAS_I_1_C_1 : begin
        fsm_output = 92'b1000000000000000000000000000000000000000000;
        state_var_NS = BIAS_I_1_C_2;
      end
      BIAS_I_1_C_2 : begin
        fsm_output = 92'b10000000000000000000000000000000000000000000;
        if ( BIAS_I_1_C_2_tr0 ) begin
          state_var_NS = BIAS_J_1_C_0;
        end
        else begin
          state_var_NS = BIAS_I_1_C_0;
        end
      end
      BIAS_J_1_C_0 : begin
        fsm_output = 92'b100000000000000000000000000000000000000000000;
        if ( BIAS_J_1_C_0_tr0 ) begin
          state_var_NS = FOR_L_1_C_0;
        end
        else begin
          state_var_NS = BIAS_I_1_C_0;
        end
      end
      FOR_L_1_C_0 : begin
        fsm_output = 92'b1000000000000000000000000000000000000000000000;
        if ( FOR_L_1_C_0_tr0 ) begin
          state_var_NS = FOR_J_3_C_0;
        end
        else begin
          state_var_NS = FOR_B_2_C_0;
        end
      end
      FOR_J_3_C_0 : begin
        fsm_output = 92'b10000000000000000000000000000000000000000000000;
        state_var_NS = FOR_I_3_C_0;
      end
      FOR_I_3_C_0 : begin
        fsm_output = 92'b100000000000000000000000000000000000000000000000;
        state_var_NS = FOR_A_3_C_0;
      end
      FOR_A_3_C_0 : begin
        fsm_output = 92'b1000000000000000000000000000000000000000000000000;
        state_var_NS = FOR_A_3_C_1;
      end
      FOR_A_3_C_1 : begin
        fsm_output = 92'b10000000000000000000000000000000000000000000000000;
        if ( FOR_A_3_C_1_tr0 ) begin
          state_var_NS = FOR_B_3_C_0;
        end
        else begin
          state_var_NS = FOR_A_3_C_0;
        end
      end
      FOR_B_3_C_0 : begin
        fsm_output = 92'b100000000000000000000000000000000000000000000000000;
        state_var_NS = FOR_B_3_C_1;
      end
      FOR_B_3_C_1 : begin
        fsm_output = 92'b1000000000000000000000000000000000000000000000000000;
        if ( FOR_B_3_C_1_tr0 ) begin
          state_var_NS = FOR_I_3_C_1;
        end
        else begin
          state_var_NS = FOR_A_3_C_0;
        end
      end
      FOR_I_3_C_1 : begin
        fsm_output = 92'b10000000000000000000000000000000000000000000000000000;
        if ( FOR_I_3_C_1_tr0 ) begin
          state_var_NS = FOR_J_3_C_1;
        end
        else begin
          state_var_NS = FOR_I_3_C_0;
        end
      end
      FOR_J_3_C_1 : begin
        fsm_output = 92'b100000000000000000000000000000000000000000000000000000;
        if ( FOR_J_3_C_1_tr0 ) begin
          state_var_NS = FOR_K_3_C_0;
        end
        else begin
          state_var_NS = FOR_J_3_C_0;
        end
      end
      FOR_K_3_C_0 : begin
        fsm_output = 92'b1000000000000000000000000000000000000000000000000000000;
        if ( FOR_K_3_C_0_tr0 ) begin
          state_var_NS = INIT_I_2_C_0;
        end
        else begin
          state_var_NS = FOR_J_3_C_0;
        end
      end
      INIT_I_2_C_0 : begin
        fsm_output = 92'b10000000000000000000000000000000000000000000000000000000;
        state_var_NS = INIT_I_2_C_1;
      end
      INIT_I_2_C_1 : begin
        fsm_output = 92'b100000000000000000000000000000000000000000000000000000000;
        if ( INIT_I_2_C_1_tr0 ) begin
          state_var_NS = INIT_J_2_C_0;
        end
        else begin
          state_var_NS = INIT_I_2_C_0;
        end
      end
      INIT_J_2_C_0 : begin
        fsm_output = 92'b1000000000000000000000000000000000000000000000000000000000;
        if ( INIT_J_2_C_0_tr0 ) begin
          state_var_NS = INIT_L_2_C_0;
        end
        else begin
          state_var_NS = INIT_I_2_C_0;
        end
      end
      INIT_L_2_C_0 : begin
        fsm_output = 92'b10000000000000000000000000000000000000000000000000000000000;
        if ( INIT_L_2_C_0_tr0 ) begin
          state_var_NS = FOR_B_4_C_0;
        end
        else begin
          state_var_NS = INIT_I_2_C_0;
        end
      end
      FOR_B_4_C_0 : begin
        fsm_output = 92'b100000000000000000000000000000000000000000000000000000000000;
        state_var_NS = FOR_B_4_C_1;
      end
      FOR_B_4_C_1 : begin
        fsm_output = 92'b1000000000000000000000000000000000000000000000000000000000000;
        if ( FOR_B_4_C_1_tr0 ) begin
          state_var_NS = FOR_A_4_C_0;
        end
        else begin
          state_var_NS = FOR_B_4_C_0;
        end
      end
      FOR_A_4_C_0 : begin
        fsm_output = 92'b10000000000000000000000000000000000000000000000000000000000000;
        if ( FOR_A_4_C_0_tr0 ) begin
          state_var_NS = FOR_I_4_C_0;
        end
        else begin
          state_var_NS = FOR_B_4_C_0;
        end
      end
      FOR_I_4_C_0 : begin
        fsm_output = 92'b100000000000000000000000000000000000000000000000000000000000000;
        state_var_NS = FOR_I_4_C_1;
      end
      FOR_I_4_C_1 : begin
        fsm_output = 92'b1000000000000000000000000000000000000000000000000000000000000000;
        state_var_NS = FOR_I_4_C_2;
      end
      FOR_I_4_C_2 : begin
        fsm_output = 92'b10000000000000000000000000000000000000000000000000000000000000000;
        if ( FOR_I_4_C_2_tr0 ) begin
          state_var_NS = FOR_J_4_C_0;
        end
        else begin
          state_var_NS = FOR_B_4_C_0;
        end
      end
      FOR_J_4_C_0 : begin
        fsm_output = 92'b100000000000000000000000000000000000000000000000000000000000000000;
        if ( FOR_J_4_C_0_tr0 ) begin
          state_var_NS = FOR_K_4_C_0;
        end
        else begin
          state_var_NS = FOR_B_4_C_0;
        end
      end
      FOR_K_4_C_0 : begin
        fsm_output = 92'b1000000000000000000000000000000000000000000000000000000000000000000;
        if ( FOR_K_4_C_0_tr0 ) begin
          state_var_NS = BIAS_I_2_C_0;
        end
        else begin
          state_var_NS = FOR_B_4_C_0;
        end
      end
      BIAS_I_2_C_0 : begin
        fsm_output = 92'b10000000000000000000000000000000000000000000000000000000000000000000;
        state_var_NS = BIAS_I_2_C_1;
      end
      BIAS_I_2_C_1 : begin
        fsm_output = 92'b100000000000000000000000000000000000000000000000000000000000000000000;
        state_var_NS = BIAS_I_2_C_2;
      end
      BIAS_I_2_C_2 : begin
        fsm_output = 92'b1000000000000000000000000000000000000000000000000000000000000000000000;
        if ( BIAS_I_2_C_2_tr0 ) begin
          state_var_NS = BIAS_J_2_C_0;
        end
        else begin
          state_var_NS = BIAS_I_2_C_0;
        end
      end
      BIAS_J_2_C_0 : begin
        fsm_output = 92'b10000000000000000000000000000000000000000000000000000000000000000000000;
        if ( BIAS_J_2_C_0_tr0 ) begin
          state_var_NS = FOR_L_2_C_0;
        end
        else begin
          state_var_NS = BIAS_I_2_C_0;
        end
      end
      FOR_L_2_C_0 : begin
        fsm_output = 92'b100000000000000000000000000000000000000000000000000000000000000000000000;
        if ( FOR_L_2_C_0_tr0 ) begin
          state_var_NS = FOR_J_5_C_0;
        end
        else begin
          state_var_NS = FOR_B_4_C_0;
        end
      end
      FOR_J_5_C_0 : begin
        fsm_output = 92'b1000000000000000000000000000000000000000000000000000000000000000000000000;
        state_var_NS = FOR_I_5_C_0;
      end
      FOR_I_5_C_0 : begin
        fsm_output = 92'b10000000000000000000000000000000000000000000000000000000000000000000000000;
        state_var_NS = FOR_A_5_C_0;
      end
      FOR_A_5_C_0 : begin
        fsm_output = 92'b100000000000000000000000000000000000000000000000000000000000000000000000000;
        state_var_NS = FOR_A_5_C_1;
      end
      FOR_A_5_C_1 : begin
        fsm_output = 92'b1000000000000000000000000000000000000000000000000000000000000000000000000000;
        if ( FOR_A_5_C_1_tr0 ) begin
          state_var_NS = FOR_B_5_C_0;
        end
        else begin
          state_var_NS = FOR_A_5_C_0;
        end
      end
      FOR_B_5_C_0 : begin
        fsm_output = 92'b10000000000000000000000000000000000000000000000000000000000000000000000000000;
        state_var_NS = FOR_B_5_C_1;
      end
      FOR_B_5_C_1 : begin
        fsm_output = 92'b100000000000000000000000000000000000000000000000000000000000000000000000000000;
        if ( FOR_B_5_C_1_tr0 ) begin
          state_var_NS = FOR_I_5_C_1;
        end
        else begin
          state_var_NS = FOR_A_5_C_0;
        end
      end
      FOR_I_5_C_1 : begin
        fsm_output = 92'b1000000000000000000000000000000000000000000000000000000000000000000000000000000;
        if ( FOR_I_5_C_1_tr0 ) begin
          state_var_NS = FOR_J_5_C_1;
        end
        else begin
          state_var_NS = FOR_I_5_C_0;
        end
      end
      FOR_J_5_C_1 : begin
        fsm_output = 92'b10000000000000000000000000000000000000000000000000000000000000000000000000000000;
        if ( FOR_J_5_C_1_tr0 ) begin
          state_var_NS = FOR_K_5_C_0;
        end
        else begin
          state_var_NS = FOR_J_5_C_0;
        end
      end
      FOR_K_5_C_0 : begin
        fsm_output = 92'b100000000000000000000000000000000000000000000000000000000000000000000000000000000;
        if ( FOR_K_5_C_0_tr0 ) begin
          state_var_NS = FOR_K_6_C_0;
        end
        else begin
          state_var_NS = FOR_J_5_C_0;
        end
      end
      FOR_K_6_C_0 : begin
        fsm_output = 92'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        state_var_NS = FOR_K_6_C_1;
      end
      FOR_K_6_C_1 : begin
        fsm_output = 92'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        state_var_NS = FOR_K_6_C_2;
      end
      FOR_K_6_C_2 : begin
        fsm_output = 92'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        if ( FOR_K_6_C_2_tr0 ) begin
          state_var_NS = FOR_J_6_C_0;
        end
        else begin
          state_var_NS = FOR_K_6_C_0;
        end
      end
      FOR_J_6_C_0 : begin
        fsm_output = 92'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        if ( FOR_J_6_C_0_tr0 ) begin
          state_var_NS = FOR_I_6_C_0;
        end
        else begin
          state_var_NS = FOR_K_6_C_0;
        end
      end
      FOR_I_6_C_0 : begin
        fsm_output = 92'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        if ( FOR_I_6_C_0_tr0 ) begin
          state_var_NS = FOR_J_7_C_0;
        end
        else begin
          state_var_NS = FOR_K_6_C_0;
        end
      end
      FOR_J_7_C_0 : begin
        fsm_output = 92'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        state_var_NS = FOR_K_7_C_0;
      end
      FOR_K_7_C_0 : begin
        fsm_output = 92'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        state_var_NS = FOR_K_7_C_1;
      end
      FOR_K_7_C_1 : begin
        fsm_output = 92'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        if ( FOR_K_7_C_1_tr0 ) begin
          state_var_NS = FOR_J_7_C_1;
        end
        else begin
          state_var_NS = FOR_K_7_C_0;
        end
      end
      FOR_J_7_C_1 : begin
        fsm_output = 92'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        if ( FOR_J_7_C_1_tr0 ) begin
          state_var_NS = for_C_0;
        end
        else begin
          state_var_NS = FOR_J_7_C_0;
        end
      end
      for_C_0 : begin
        fsm_output = 92'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        if ( for_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = for_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 92'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 92'b1;
        state_var_NS = core_rlp_C_1;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= core_rlp_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    CNN_main_simple_core
// ------------------------------------------------------------------


module CNN_main_simple_core (
  clk, rst, image_rsc_triosy_lz, F_1_rsc_triosy_lz, B_1_rsc_triosy_lz, F_2_rsc_triosy_lz,
      B_2_rsc_triosy_lz, F_3_rsc_triosy_lz, B_3_rsc_triosy_lz, P_W_rsc_triosy_lz,
      P_B_rsc_triosy_lz, index_rsc_dat, index_rsc_triosy_lz, image_rsci_radr_d, image_rsci_q_d,
      F_1_rsci_radr_d, F_1_rsci_q_d, B_1_rsci_radr_d, B_1_rsci_re_d, B_1_rsci_q_d,
      F_2_rsci_radr_d, F_2_rsci_re_d, F_2_rsci_q_d, B_2_rsci_radr_d, B_2_rsci_re_d,
      B_2_rsci_q_d, F_3_rsci_radr_d, F_3_rsci_re_d, F_3_rsci_q_d, B_3_rsci_radr_d,
      B_3_rsci_re_d, B_3_rsci_q_d, P_W_rsci_radr_d, P_W_rsci_re_d, P_W_rsci_q_d,
      P_B_rsci_radr_d, P_B_rsci_re_d, P_B_rsci_q_d, memory_1_rsci_radr_d, memory_1_rsci_wadr_d,
      memory_1_rsci_d_d, memory_1_rsci_we_d, memory_1_rsci_re_d, memory_1_rsci_q_d,
      memory_2_rsci_radr_d, memory_2_rsci_wadr_d, memory_2_rsci_d_d, memory_2_rsci_we_d,
      memory_2_rsci_re_d, memory_2_rsci_q_d, image_rsci_re_d_pff
);
  input clk;
  input rst;
  output image_rsc_triosy_lz;
  output F_1_rsc_triosy_lz;
  output B_1_rsc_triosy_lz;
  output F_2_rsc_triosy_lz;
  output B_2_rsc_triosy_lz;
  output F_3_rsc_triosy_lz;
  output B_3_rsc_triosy_lz;
  output P_W_rsc_triosy_lz;
  output P_B_rsc_triosy_lz;
  output [3:0] index_rsc_dat;
  output index_rsc_triosy_lz;
  output [10:0] image_rsci_radr_d;
  input [15:0] image_rsci_q_d;
  output [10:0] F_1_rsci_radr_d;
  input [15:0] F_1_rsci_q_d;
  output [5:0] B_1_rsci_radr_d;
  output B_1_rsci_re_d;
  input [15:0] B_1_rsci_q_d;
  output [14:0] F_2_rsci_radr_d;
  output F_2_rsci_re_d;
  input [15:0] F_2_rsci_q_d;
  output [4:0] B_2_rsci_radr_d;
  output B_2_rsci_re_d;
  input [15:0] B_2_rsci_q_d;
  output [12:0] F_3_rsci_radr_d;
  output F_3_rsci_re_d;
  input [15:0] F_3_rsci_q_d;
  output [4:0] B_3_rsci_radr_d;
  output B_3_rsci_re_d;
  input [15:0] B_3_rsci_q_d;
  output [10:0] P_W_rsci_radr_d;
  output P_W_rsci_re_d;
  input [15:0] P_W_rsci_q_d;
  output [3:0] P_B_rsci_radr_d;
  output P_B_rsci_re_d;
  input [15:0] P_B_rsci_q_d;
  output [10:0] memory_1_rsci_radr_d;
  output [10:0] memory_1_rsci_wadr_d;
  output [15:0] memory_1_rsci_d_d;
  output memory_1_rsci_we_d;
  output memory_1_rsci_re_d;
  input [15:0] memory_1_rsci_q_d;
  output [10:0] memory_2_rsci_radr_d;
  output [10:0] memory_2_rsci_wadr_d;
  output [15:0] memory_2_rsci_d_d;
  output memory_2_rsci_we_d;
  output memory_2_rsci_re_d;
  input [15:0] memory_2_rsci_q_d;
  output image_rsci_re_d_pff;


  // Interconnect Declarations
  reg [3:0] index_rsci_idat;
  wire [91:0] fsm_output;
  wire or_dcpl_53;
  wire and_dcpl_6;
  wire and_dcpl_133;
  wire or_dcpl_130;
  wire or_dcpl_131;
  wire and_dcpl_136;
  wire or_dcpl_134;
  wire or_dcpl_135;
  wire and_dcpl_141;
  wire or_dcpl_139;
  wire or_dcpl_140;
  wire or_dcpl_142;
  wire or_tmp_111;
  wire or_tmp_117;
  wire or_tmp_125;
  wire or_tmp_376;
  wire or_tmp_379;
  wire or_tmp_380;
  wire or_tmp_383;
  wire or_tmp_392;
  wire or_tmp_393;
  wire or_tmp_405;
  wire or_tmp_406;
  wire or_tmp_418;
  wire or_tmp_419;
  wire or_tmp_431;
  wire or_tmp_432;
  wire or_tmp_444;
  wire or_tmp_445;
  wire or_tmp_457;
  wire or_tmp_458;
  wire or_tmp_470;
  wire or_tmp_471;
  wire or_tmp_483;
  wire or_tmp_484;
  wire or_tmp_496;
  wire or_tmp_497;
  wire FOR_B_4_oelse_acc_tmp_15;
  wire FOR_B_2_oelse_acc_tmp_14;
  wire FOR_B_oelse_acc_tmp_13;
  wire and_4_cse;
  wire and_10_cse;
  wire and_16_cse;
  wire and_285_cse;
  wire and_283_cse;
  wire and_316_cse;
  wire and_318_cse;
  wire and_317_cse;
  wire and_386_cse;
  wire and_307_cse;
  reg FOR_K_7_slc_FOR_K_7_acc_6_itm;
  reg FOR_K_7_mux_28_itm;
  reg [13:0] FOR_K_7_mux_29_itm;
  reg FOR_K_7_mux_30_itm;
  wire FOR_J_7_and_stg_2_1_sva_1;
  wire FOR_J_7_and_stg_2_0_sva_1;
  wire FOR_J_7_and_stg_1_3_sva_1;
  wire FOR_J_7_and_stg_1_2_sva_1;
  wire FOR_J_7_and_stg_1_1_sva_1;
  wire FOR_J_7_and_stg_1_0_sva_1;
  reg FOR_K_6_slc_FOR_K_6_acc_3_itm;
  reg [1:0] MP3_simple_a_1_0_sva;
  reg BIAS_I_2_slc_BIAS_I_2_acc_2_itm;
  reg [14:0] BIAS_I_2_slc_15_1_itm;
  reg FOR_I_4_slc_FOR_I_4_acc_2_itm;
  reg CR3_simple_aux_15_lpi_7_dfm;
  reg [13:0] CR3_simple_aux_14_1_lpi_7_dfm;
  reg CR3_simple_aux_0_lpi_7_dfm;
  reg CR3_simple_aux_15_lpi_7;
  reg [13:0] CR3_simple_aux_14_1_lpi_7;
  reg CR3_simple_aux_0_lpi_7;
  reg BIAS_I_1_slc_BIAS_I_1_acc_2_itm;
  reg [14:0] BIAS_I_1_slc_15_1_itm;
  reg FOR_I_2_slc_FOR_I_2_acc_2_itm;
  reg CR2_simple_aux_15_lpi_7_dfm;
  reg [13:0] CR2_simple_aux_14_1_lpi_7_dfm;
  reg CR2_simple_aux_0_lpi_7_dfm;
  reg CR2_simple_aux_15_lpi_7;
  reg [13:0] CR2_simple_aux_14_1_lpi_7;
  reg CR2_simple_aux_0_lpi_7;
  reg BIAS_I_slc_BIAS_I_acc_2_itm;
  reg [14:0] BIAS_I_slc_15_1_itm;
  reg FOR_I_slc_FOR_I_acc_2_itm;
  reg CR1_simple_aux_15_lpi_7_dfm;
  reg [13:0] CR1_simple_aux_14_1_lpi_7_dfm;
  reg CR1_simple_aux_0_lpi_7_dfm;
  reg CR1_simple_aux_15_lpi_7;
  reg [13:0] CR1_simple_aux_14_1_lpi_7;
  reg CR1_simple_aux_0_lpi_7;
  reg FOR_J_7_and_21_cse_sva;
  reg FOR_J_7_and_20_cse_sva;
  reg FOR_J_7_and_19_cse_sva;
  reg FOR_J_7_and_18_cse_sva;
  reg FOR_J_7_and_17_cse_sva;
  reg FOR_J_7_and_16_cse_sva;
  reg FOR_J_7_and_15_cse_sva;
  reg FOR_J_7_and_14_cse_sva;
  reg FOR_J_7_and_13_cse_sva;
  reg FOR_J_7_and_12_cse_sva;
  reg [3:0] perceptron_simple_j_3_0_sva;
  reg max_sva_15;
  reg [13:0] max_sva_14_1;
  reg max_sva_0;
  wire for_slc_Prob_16_15_0_cse_sva_15_1;
  wire [13:0] for_slc_Prob_16_15_0_cse_sva_14_1_1;
  wire for_slc_Prob_16_15_0_cse_sva_0_1;
  reg [15:0] MP3_simple_bigger_lpi_6;
  reg [15:0] MP2_simple_bigger_lpi_6;
  reg [15:0] MP1_simple_bigger_lpi_6;
  reg [1:0] CR1_simple_b_1_0_sva_1;
  wire [16:0] FOR_K_7_acc_7_psp_sva_1;
  wire [17:0] nl_FOR_K_7_acc_7_psp_sva_1;
  wire [18:0] FOR_B_if_acc_psp_sva_1;
  wire [19:0] nl_FOR_B_if_acc_psp_sva_1;
  wire [4:0] FOR_A_1_if_asn_MP1_simple_add_M_10_FOR_A_1_if_acc_sdt;
  wire [5:0] nl_FOR_A_1_if_asn_MP1_simple_add_M_10_FOR_A_1_if_acc_sdt;
  wire [4:0] INIT_I_asn_CR1_simple_add_AF_10_INIT_I_acc_sdt;
  wire [5:0] nl_INIT_I_asn_CR1_simple_add_AF_10_INIT_I_acc_sdt;
  wire or_220_ssc;
  wire [4:0] FOR_B_4_if_acc_10_sdt_4_0_1;
  wire [5:0] nl_FOR_B_4_if_acc_10_sdt_4_0_1;
  reg reg_index_rsc_triosy_obj_ld_cse;
  wire reg_CR1_simple_CR1_simple_aux_or_1_cse;
  wire or_125_cse;
  wire reg_CR2_simple_CR2_simple_aux_or_1_cse;
  wire reg_CR3_simple_CR3_simple_aux_or_1_cse;
  wire FOR_B_2_if_FOR_B_2_if_or_cse;
  wire or_332_cse;
  wire or_400_cse;
  wire or_468_cse;
  wire FOR_B_4_if_FOR_B_4_if_or_cse;
  wire reg_CR1_simple_l_1_6_0_sva_5_CR1_simple_l_or_cse;
  wire reg_MP3_simple_b_1_MP3_simple_b_or_cse;
  wire memory_1_nor_1_seb;
  wire memory_1_or_1_seb;
  wire memory_1_or_seb;
  wire [7:0] FOR_K_7_acc_8_sdt_1;
  wire [8:0] nl_FOR_K_7_acc_8_sdt_1;
  reg [7:0] perceptron_simple_k_7_0_sva;
  reg [4:0] CR3_simple_l_4_0_sva;
  reg [1:0] CR2_simple_a_1_0_sva;
  reg [5:0] CR2_simple_k_6_0_sva_5_0_1;
  reg [4:0] CR2_simple_l_5_0_sva_4_0_1;
  reg [5:0] CR1_simple_l_6_0_sva_5_0_1;
  reg [1:0] CR1_simple_k_1_0_sva;
  wire [6:0] FOR_B_if_acc_10_psp_1;
  wire [7:0] nl_FOR_B_if_acc_10_psp_1;
  wire [5:0] FOR_B_if_acc_5_sdt_1;
  wire [6:0] nl_FOR_B_if_acc_5_sdt_1;
  wire [6:0] FOR_B_2_if_acc_8_sdt_1;
  wire [7:0] nl_FOR_B_2_if_acc_8_sdt_1;
  wire [5:0] FOR_B_2_if_acc_9_psp_1;
  wire [6:0] nl_FOR_B_2_if_acc_9_psp_1;
  wire [6:0] FOR_B_4_if_acc_11_sdt_1;
  wire [7:0] nl_FOR_B_4_if_acc_11_sdt_1;
  reg [4:0] CR3_simple_k_5_0_sva_4_0;
  reg [4:0] reshape_simple_k_4_0_sva;
  wire memory_2_rsci_radr_d_mx0c0;
  wire [4:0] CR2_simple_j_aux_4_0_sva_1;
  wire [5:0] nl_CR2_simple_j_aux_4_0_sva_1;
  wire [4:0] FOR_B_4_if_acc_6_sdt_1;
  wire [5:0] nl_FOR_B_4_if_acc_6_sdt_1;
  wire [3:0] CR3_simple_j_aux_3_0_sva_1;
  wire [4:0] nl_CR3_simple_j_aux_3_0_sva_1;
  wire [6:0] FOR_B_1_if_acc_3_sdt_1;
  wire [7:0] nl_FOR_B_1_if_acc_3_sdt_1;
  reg [5:0] MP1_simple_k_6_0_sva_5_0;
  reg [4:0] MP2_simple_k_5_0_sva_4_0;
  reg [4:0] MP3_simple_k_4_0_sva;
  wire memory_2_rsci_wadr_d_mx0c0;
  reg [3:0] MP1_simple_i_N_3_0_sva_1;
  wire [2:0] FOR_B_3_if_acc_sdt_1;
  wire [3:0] nl_FOR_B_3_if_acc_sdt_1;
  reg [2:0] MP2_simple_i_N_2_0_sva_1;
  reg [1:0] CR3_simple_a_1_0_sva;
  reg [1:0] CR1_simple_a_1_0_sva;
  reg [15:0] MP1_simple_bigger_lpi_6_dfm_1;
  reg [15:0] MP2_simple_bigger_lpi_6_dfm_1;
  reg [15:0] MP3_simple_bigger_lpi_6_dfm_1;
  reg [4:0] CR1_simple_j_2_4_0_sva;
  reg [4:0] CR1_simple_j_4_0_sva;
  wire [3:0] FOR_A_1_oelse_acc_1_ncse_sva_2;
  wire [4:0] nl_FOR_A_1_oelse_acc_1_ncse_sva_2;
  reg [3:0] CR2_simple_j_2_3_0_sva;
  reg [3:0] CR2_simple_j_3_0_sva;
  wire [2:0] FOR_A_3_oelse_acc_1_ncse_sva_2;
  wire [3:0] nl_FOR_A_3_oelse_acc_1_ncse_sva_2;
  reg [1:0] MP1_simple_a_1_0_sva;
  reg [1:0] MP2_simple_a_1_0_sva;
  reg [2:0] CR3_simple_j_2_2_0_sva;
  reg [2:0] CR3_simple_j_2_0_sva;
  reg [10:0] reshape_simple_add_N_10_0_lpi_4;
  wire [4:0] INIT_I_2_acc_6_sdt_1;
  wire [5:0] nl_INIT_I_2_acc_6_sdt_1;
  reg [4:0] CR3_simple_l_1_4_0_sva;
  reg [4:0] CR1_simple_j_1_4_0_sva;
  reg [3:0] CR2_simple_j_1_3_0_sva;
  reg [2:0] CR3_simple_j_1_2_0_sva;
  wire [2:0] z_out;
  wire [2:0] z_out_2;
  wire [3:0] nl_z_out_2;
  wire [2:0] z_out_3;
  wire [3:0] nl_z_out_3;
  wire [2:0] z_out_4;
  wire [3:0] z_out_5;
  wire [4:0] nl_z_out_5;
  wire [2:0] z_out_6;
  wire [3:0] nl_z_out_6;
  wire [3:0] z_out_7;
  wire [4:0] nl_z_out_7;
  wire [3:0] z_out_8;
  wire [4:0] nl_z_out_8;
  wire [4:0] z_out_9;
  wire [5:0] nl_z_out_9;
  wire [5:0] z_out_10;
  wire [6:0] nl_z_out_10;
  wire [5:0] z_out_11;
  wire [6:0] nl_z_out_11;
  wire [4:0] z_out_12;
  wire [5:0] nl_z_out_12;
  wire [6:0] z_out_13;
  wire [7:0] nl_z_out_13;
  wire [5:0] z_out_16;
  wire [6:0] nl_z_out_16;
  wire [1:0] z_out_17;
  wire [2:0] nl_z_out_17;
  wire [4:0] z_out_19;
  wire [5:0] nl_z_out_19;
  wire [4:0] z_out_20;
  wire [5:0] nl_z_out_20;
  wire [4:0] z_out_21;
  wire [5:0] nl_z_out_21;
  wire [16:0] z_out_22;
  wire [4:0] z_out_23;
  wire [5:0] nl_z_out_23;
  wire [19:0] z_out_24;
  wire [20:0] nl_z_out_24;
  wire [3:0] z_out_25;
  wire [4:0] nl_z_out_25;
  wire [3:0] z_out_26;
  wire [4:0] nl_z_out_26;
  reg [4:0] CR1_simple_i_1_4_0_sva;
  reg [4:0] CR1_simple_i_1_4_0_sva_1;
  reg [4:0] CR1_simple_i_2_4_0_sva;
  reg [1:0] CR1_simple_b_1_0_sva;
  reg [4:0] CR1_simple_i_2_4_0_sva_1;
  reg [4:0] CR1_simple_i_4_0_sva;
  reg [4:0] CR1_simple_i_4_0_sva_1;
  reg [3:0] MP1_simple_j_N_3_0_sva;
  reg [3:0] MP1_simple_j_4_1_sva;
  reg [3:0] MP1_simple_j_N_3_0_sva_1;
  reg [3:0] MP1_simple_i_N_3_0_sva;
  reg [3:0] MP1_simple_i_4_1_sva;
  reg [1:0] MP1_simple_b_1_0_sva;
  reg [3:0] CR2_simple_i_1_3_0_sva;
  reg [3:0] CR2_simple_i_1_3_0_sva_1;
  reg [3:0] CR2_simple_i_2_3_0_sva;
  reg [1:0] CR2_simple_b_1_0_sva;
  reg [3:0] CR2_simple_i_2_3_0_sva_1;
  reg [3:0] CR2_simple_i_3_0_sva;
  reg [3:0] CR2_simple_i_3_0_sva_1;
  reg [2:0] MP2_simple_j_N_2_0_sva;
  reg [2:0] MP2_simple_j_3_1_sva;
  reg [2:0] MP2_simple_j_N_2_0_sva_1;
  reg [2:0] MP2_simple_i_N_2_0_sva;
  reg [2:0] MP2_simple_i_3_1_sva;
  reg [1:0] MP2_simple_b_1_0_sva;
  reg [2:0] CR3_simple_i_1_2_0_sva;
  reg [2:0] CR3_simple_i_1_2_0_sva_1;
  reg [2:0] CR3_simple_i_2_2_0_sva;
  reg [1:0] CR3_simple_b_1_0_sva;
  reg [2:0] CR3_simple_i_2_2_0_sva_1;
  reg [2:0] CR3_simple_i_2_0_sva;
  reg [2:0] CR3_simple_i_2_0_sva_1;
  reg [1:0] MP3_simple_j_2_1_sva;
  reg [1:0] MP3_simple_j_N_1_0_sva_1;
  reg [1:0] MP3_simple_i_2_1_sva;
  reg [1:0] MP3_simple_i_N_1_0_sva_1;
  reg [1:0] MP3_simple_b_1_0_sva;
  reg [1:0] reshape_simple_i_1_0_sva;
  reg [1:0] reshape_simple_j_1_0_sva;
  reg [10:0] reshape_simple_add_N_10_0_sva_1;
  wire [11:0] nl_reshape_simple_add_N_10_0_sva_1;
  reg [4:0] reshape_simple_k_4_0_sva_1;
  reg [13:0] Prob_4_14_1_sva_1;
  reg Prob_4_0_sva_1;
  reg Prob_4_15_sva_1;
  reg [13:0] Prob_5_14_1_sva_1;
  reg Prob_5_0_sva_1;
  reg Prob_5_15_sva_1;
  reg [13:0] Prob_3_14_1_sva_1;
  reg Prob_3_0_sva_1;
  reg Prob_3_15_sva_1;
  reg [13:0] Prob_6_14_1_sva_1;
  reg Prob_6_0_sva_1;
  reg Prob_6_15_sva_1;
  reg [13:0] Prob_2_14_1_sva_1;
  reg Prob_2_0_sva_1;
  reg Prob_2_15_sva_1;
  reg [13:0] Prob_7_14_1_sva_1;
  reg Prob_7_0_sva_1;
  reg Prob_7_15_sva_1;
  reg [13:0] Prob_1_14_1_sva_1;
  reg Prob_1_0_sva_1;
  reg Prob_1_15_sva_1;
  reg [13:0] Prob_8_14_1_sva_1;
  reg Prob_8_0_sva_1;
  reg Prob_8_15_sva_1;
  reg [13:0] Prob_9_14_1_sva_1;
  reg Prob_9_0_sva_1;
  reg Prob_9_15_sva_1;
  reg [13:0] Prob_4_14_1_sva_2;
  reg Prob_4_0_sva_2;
  reg Prob_4_15_sva_2;
  reg [13:0] Prob_5_14_1_sva_2;
  reg Prob_5_0_sva_2;
  reg Prob_5_15_sva_2;
  reg [13:0] Prob_3_14_1_sva_2;
  reg Prob_3_0_sva_2;
  reg Prob_3_15_sva_2;
  reg [13:0] Prob_6_14_1_sva_2;
  reg Prob_6_0_sva_2;
  reg Prob_6_15_sva_2;
  reg [13:0] Prob_2_14_1_sva_2;
  reg Prob_2_0_sva_2;
  reg Prob_2_15_sva_2;
  reg [13:0] Prob_7_14_1_sva_2;
  reg Prob_7_0_sva_2;
  reg Prob_7_15_sva_2;
  reg [13:0] Prob_1_14_1_sva_2;
  reg Prob_1_0_sva_2;
  reg Prob_1_15_sva_2;
  reg [13:0] Prob_8_14_1_sva_2;
  reg Prob_8_0_sva_2;
  reg Prob_8_15_sva_2;
  reg [13:0] Prob_9_14_1_sva_2;
  reg Prob_9_0_sva_2;
  reg Prob_9_15_sva_2;
  reg [7:0] perceptron_simple_k_7_0_sva_1;
  reg [3:0] k_sva;
  reg FOR_B_lor_2_lpi_7_dfm_st;
  reg FOR_B_2_lor_2_lpi_7_dfm_st;
  reg FOR_B_4_lor_2_lpi_7_dfm_st;
  reg [5:0] CR1_simple_l_1_6_0_sva_5_0;
  reg [4:0] CR2_simple_l_1_5_0_sva_4_0;
  reg Prob_0_sva_1_15;
  reg [13:0] Prob_0_sva_1_14_1;
  reg Prob_0_sva_1_0;
  reg Prob_0_sva_2_15;
  reg [13:0] Prob_0_sva_2_14_1;
  reg Prob_0_sva_2_0;
  reg MP3_simple_j_N_1_0_sva_1_1;
  reg MP3_simple_j_N_1_0_sva_0;
  reg MP3_simple_i_N_1_0_sva_1_1;
  reg MP3_simple_i_N_1_0_sva_0;
  wire CR1_simple_aux_15_lpi_7_mx1;
  wire [13:0] CR1_simple_aux_14_1_lpi_7_mx1;
  wire CR1_simple_aux_0_lpi_7_mx1;
  wire [5:0] FOR_B_acc_1_psp_sva_1;
  wire [6:0] nl_FOR_B_acc_1_psp_sva_1;
  wire FOR_B_if_nor_ovfl_sva_1;
  wire FOR_B_if_and_unfl_sva_1;
  wire [15:0] MP1_simple_bigger_lpi_6_mx1;
  wire CR2_simple_aux_15_lpi_7_mx1;
  wire [13:0] CR2_simple_aux_14_1_lpi_7_mx1;
  wire CR2_simple_aux_0_lpi_7_mx1;
  wire [4:0] FOR_B_2_acc_1_psp_sva_1;
  wire [5:0] nl_FOR_B_2_acc_1_psp_sva_1;
  wire FOR_B_2_if_nor_ovfl_sva_1;
  wire FOR_B_2_if_and_unfl_sva_1;
  wire [15:0] MP2_simple_bigger_lpi_6_mx1;
  wire CR3_simple_aux_15_lpi_7_mx1;
  wire [13:0] CR3_simple_aux_14_1_lpi_7_mx1;
  wire CR3_simple_aux_0_lpi_7_mx1;
  wire [3:0] FOR_B_4_acc_1_psp_1_sva_1;
  wire [4:0] nl_FOR_B_4_acc_1_psp_1_sva_1;
  wire [15:0] MP3_simple_bigger_lpi_6_mx1;
  wire reshape_simple_add_N_10_0_lpi_4_mx0c1;
  wire [7:0] perceptron_simple_k_7_0_sva_2;
  wire [8:0] nl_perceptron_simple_k_7_0_sva_2;
  wire FOR_K_7_FOR_K_7_nor_2_psp_sva_1;
  wire [13:0] FOR_K_7_FOR_K_7_nor_1_psp_sva_1;
  wire FOR_K_7_nor_ovfl_sva_1;
  wire FOR_K_7_and_unfl_sva_1;
  wire [13:0] max_sva_14_1_mx1;
  wire FOR_B_oelse_2_acc_itm_13;
  wire FOR_B_2_oelse_2_acc_itm_14;
  wire [3:0] FOR_A_1_if_mux1h_4_cse;
  wire FOR_J_7_or_29_rgt;
  wire FOR_J_7_and_81_rgt;
  wire FOR_J_7_or_2_rgt;
  wire FOR_J_7_and_27_rgt;
  wire FOR_J_7_or_26_rgt;
  wire FOR_J_7_and_75_rgt;
  wire FOR_J_7_or_23_rgt;
  wire FOR_J_7_and_69_rgt;
  wire FOR_J_7_or_20_rgt;
  wire FOR_J_7_and_63_rgt;
  wire FOR_J_7_or_17_rgt;
  wire FOR_J_7_and_57_rgt;
  wire FOR_J_7_or_14_rgt;
  wire FOR_J_7_and_51_rgt;
  wire FOR_J_7_or_11_rgt;
  wire FOR_J_7_and_45_rgt;
  wire FOR_J_7_or_8_rgt;
  wire FOR_J_7_and_39_rgt;
  wire FOR_J_7_or_5_rgt;
  wire FOR_J_7_and_33_rgt;
  wire nand_cse_1;
  reg [4:0] reg_FOR_I_asn_CR1_simple_add_AF_10_FOR_I_acc_psp_cse;
  reg reg_INIT_I_slc_INIT_I_acc_2_cse;
  reg [3:0] reg_FOR_I_2_acc_11_psp_cse;
  reg [2:0] reg_FOR_I_2_acc_9_sdt_cse;
  reg reg_FOR_I_2_acc_10_psp_cse;
  reg reg_FOR_I_2_acc_8_sdt_cse;
  reg [4:0] reg_FOR_I_4_acc_11_psp_cse;
  reg [2:0] reg_FOR_I_4_acc_9_sdt_cse;
  reg reg_FOR_I_4_acc_8_sdt_2_0_cse;
  wire FOR_I_nor_2_cse;
  wire FOR_I_and_4_cse;
  wire FOR_I_6_FOR_I_6_xnor_cse;
  wire memory_1_or_2_cse;
  wire memory_1_or_5_cse;
  reg reg_FOR_A_1_lor_lpi_6_dfm_cse;
  wire [13:0] FOR_B_2_if_FOR_B_2_if_nor_cse;
  wire FOR_B_2_if_FOR_B_2_if_nor_1_cse;
  wire memory_1_or_3_cse;
  wire memory_1_or_12_cse;
  wire memory_1_or_13_cse;
  wire memory_1_or_6_cse_1;
  wire reshape_simple_add_N_or_cse;
  wire reshape_simple_add_N_or_11_cse;
  wire reshape_simple_add_N_or_2_cse;
  wire [13:0] FOR_I_nor_3_cse;
  wire FOR_I_nor_4_cse;
  wire memory_1_or_17_cse;
  wire memory_1_or_19_cse;
  wire or_141_cse;
  wire INIT_I_or_4_cse;
  wire INIT_I_or_6_cse;
  wire z_out_1_2;
  wire [1:0] z_out_14_1_0;
  wire [2:0] nl_z_out_14_1_0;
  wire [1:0] z_out_15_1_0;
  wire [2:0] nl_z_out_15_1_0;
  wire [19:0] z_out_18_31_12;
  wire [2:0] z_out_27_2_0;
  wire [3:0] nl_z_out_27_2_0;

  wire[0:0] FOR_K_7_mux_1_nl;
  wire[0:0] FOR_K_7_mux_2_nl;
  wire[0:0] Prob_Prob_nor_nl;
  wire[0:0] Prob_and_19_nl;
  wire[0:0] FOR_K_7_mux_4_nl;
  wire[0:0] FOR_K_7_mux_5_nl;
  wire[0:0] Prob_Prob_nor_1_nl;
  wire[0:0] Prob_and_17_nl;
  wire[0:0] FOR_K_7_mux_7_nl;
  wire[0:0] FOR_K_7_mux_8_nl;
  wire[0:0] Prob_Prob_nor_2_nl;
  wire[0:0] Prob_and_15_nl;
  wire[0:0] FOR_K_7_mux_10_nl;
  wire[0:0] FOR_K_7_mux_11_nl;
  wire[0:0] Prob_Prob_nor_3_nl;
  wire[0:0] Prob_and_13_nl;
  wire[0:0] FOR_K_7_mux_13_nl;
  wire[0:0] FOR_K_7_mux_14_nl;
  wire[0:0] Prob_Prob_nor_4_nl;
  wire[0:0] Prob_and_11_nl;
  wire[0:0] FOR_K_7_mux_16_nl;
  wire[0:0] FOR_K_7_mux_17_nl;
  wire[0:0] Prob_Prob_nor_5_nl;
  wire[0:0] Prob_and_9_nl;
  wire[0:0] FOR_K_7_mux_19_nl;
  wire[0:0] FOR_K_7_mux_20_nl;
  wire[0:0] Prob_Prob_nor_6_nl;
  wire[0:0] Prob_and_7_nl;
  wire[0:0] FOR_K_7_mux_22_nl;
  wire[0:0] FOR_K_7_mux_23_nl;
  wire[0:0] Prob_Prob_nor_7_nl;
  wire[0:0] Prob_and_5_nl;
  wire[0:0] FOR_K_7_mux_25_nl;
  wire[0:0] FOR_K_7_mux_26_nl;
  wire[0:0] Prob_Prob_nor_8_nl;
  wire[0:0] Prob_and_3_nl;
  wire[0:0] CR1_simple_l_not_1_nl;
  wire[0:0] CR1_simple_j_not_nl;
  wire[0:0] CR1_simple_i_nor_nl;
  wire[0:0] CR1_simple_aux_mux_14_nl;
  wire[13:0] CR1_simple_aux_mux_13_nl;
  wire[0:0] not_410_nl;
  wire[0:0] CR1_simple_aux_mux_12_nl;
  wire[0:0] not_408_nl;
  wire[0:0] MP1_simple_i_not_nl;
  wire[0:0] MP1_simple_i_N_not_nl;
  wire[0:0] MP1_simple_a_nor_nl;
  wire[0:0] MP1_simple_b_not_nl;
  wire[15:0] memory_1_mux_3_nl;
  wire[0:0] MP1_simple_bigger_not_nl;
  wire[0:0] CR1_simple_aux_mux_11_nl;
  wire[13:0] CR1_simple_aux_mux_10_nl;
  wire[0:0] not_406_nl;
  wire[0:0] CR1_simple_aux_mux_9_nl;
  wire[0:0] not_404_nl;
  wire[0:0] MP2_simple_i_not_nl;
  wire[0:0] MP2_simple_i_N_not_nl;
  wire[0:0] MP2_simple_a_nor_nl;
  wire[0:0] MP2_simple_b_not_nl;
  wire[15:0] memory_1_mux_4_nl;
  wire[0:0] MP2_simple_bigger_not_nl;
  wire[0:0] CR1_simple_aux_mux_8_nl;
  wire[13:0] CR1_simple_aux_mux_7_nl;
  wire[0:0] not_402_nl;
  wire[0:0] CR1_simple_aux_mux_6_nl;
  wire[0:0] MP3_simple_i_not_nl;
  wire[0:0] MP3_simple_a_not_nl;
  wire[0:0] MP3_simple_b_not_nl;
  wire[15:0] memory_1_mux_5_nl;
  wire[0:0] MP3_simple_bigger_not_nl;
  wire[0:0] FOR_K_7_mux_28_nl;
  wire[0:0] FOR_K_7_mux_29_nl;
  wire[0:0] Prob_Prob_nor_9_nl;
  wire[0:0] Prob_and_1_nl;
  wire[6:0] FOR_K_7_acc_nl;
  wire[7:0] nl_FOR_K_7_acc_nl;
  wire[0:0] for_mux_1_nl;
  wire[0:0] for_mux_2_nl;
  wire[13:0] FOR_B_if_FOR_B_if_nor_nl;
  wire[13:0] FOR_B_if_nor_2_nl;
  wire[0:0] FOR_B_if_FOR_B_if_nor_1_nl;
  wire[13:0] FOR_B_oelse_2_acc_nl;
  wire[14:0] nl_FOR_B_oelse_2_acc_nl;
  wire[13:0] FOR_B_oelse_acc_nl;
  wire[14:0] nl_FOR_B_oelse_acc_nl;
  wire[13:0] FOR_B_2_if_nor_2_nl;
  wire[14:0] FOR_B_2_oelse_2_acc_nl;
  wire[15:0] nl_FOR_B_2_oelse_2_acc_nl;
  wire[14:0] FOR_B_2_oelse_acc_nl;
  wire[15:0] nl_FOR_B_2_oelse_acc_nl;
  wire[4:0] FOR_B_4_if_acc_12_nl;
  wire[5:0] nl_FOR_B_4_if_acc_12_nl;
  wire[3:0] FOR_B_4_if_acc_9_nl;
  wire[4:0] nl_FOR_B_4_if_acc_9_nl;
  wire[15:0] FOR_B_4_oelse_acc_nl;
  wire[16:0] nl_FOR_B_4_oelse_acc_nl;
  wire[13:0] FOR_K_7_nor_3_nl;
  wire[4:0] BIAS_I_BIAS_I_and_2_nl;
  wire[4:0] FOR_B_if_asn_CR1_simple_add_M_10_FOR_B_if_acc_nl;
  wire[5:0] nl_FOR_B_if_asn_CR1_simple_add_M_10_FOR_B_if_acc_nl;
  wire[1:0] FOR_K_FOR_K_and_5_nl;
  wire[0:0] BIAS_I_BIAS_I_and_3_nl;
  wire[2:0] BIAS_I_2_BIAS_I_2_and_3_nl;
  wire[0:0] FOR_K_FOR_K_and_4_nl;
  wire[0:0] FOR_K_FOR_K_and_11_nl;
  wire[2:0] BIAS_I_2_BIAS_I_2_and_2_nl;
  wire[5:0] CR1_simple_l_CR1_simple_l_and_1_nl;
  wire[0:0] CR1_simple_l_nor_nl;
  wire[0:0] B_1_nor_nl;
  wire[2:0] BIAS_I_2_BIAS_I_2_and_1_nl;
  wire[0:0] BIAS_I_BIAS_I_and_1_nl;
  wire[5:0] CR2_simple_k_CR2_simple_k_and_nl;
  wire[0:0] CR2_simple_k_not_nl;
  wire[4:0] CR2_simple_l_CR2_simple_l_and_1_nl;
  wire[0:0] CR2_simple_l_not_nl;
  wire[0:0] B_2_nor_nl;
  wire[0:0] FOR_K_FOR_K_and_3_nl;
  wire[0:0] FOR_K_FOR_K_and_10_nl;
  wire[3:0] BIAS_I_1_BIAS_I_1_and_nl;
  wire[2:0] BIAS_I_2_BIAS_I_2_and_nl;
  wire[1:0] FOR_K_FOR_K_and_2_nl;
  wire[1:0] FOR_K_FOR_K_and_1_nl;
  wire[0:0] B_3_nor_nl;
  wire[7:0] FOR_K_7_FOR_K_7_and_nl;
  wire[7:0] FOR_K_7_acc_9_nl;
  wire[8:0] nl_FOR_K_7_acc_9_nl;
  wire[1:0] FOR_K_FOR_K_and_nl;
  wire[0:0] BIAS_I_BIAS_I_and_nl;
  wire[0:0] memory_1_and_1_nl;
  wire[0:0] memory_1_mux1h_1_nl;
  wire[5:0] memory_1_and_4_nl;
  wire[3:0] memory_1_mux1h_5_nl;
  wire[0:0] memory_1_mux1h_12_nl;
  wire[0:0] memory_1_mux1h_13_nl;
  wire[0:0] memory_1_and_5_nl;
  wire[0:0] memory_1_mux1h_6_nl;
  wire[0:0] memory_1_and_6_nl;
  wire[0:0] memory_1_mux1h_7_nl;
  wire[0:0] memory_1_and_7_nl;
  wire[0:0] memory_1_mux1h_8_nl;
  wire[0:0] memory_1_and_8_nl;
  wire[0:0] memory_1_mux1h_9_nl;
  wire[0:0] reshape_simple_add_N_and_nl;
  wire[0:0] reshape_simple_add_N_mux1h_nl;
  wire[5:0] reshape_simple_add_N_and_2_nl;
  wire[3:0] reshape_simple_add_N_mux1h_4_nl;
  wire[1:0] reshape_simple_add_N_mux1h_9_nl;
  wire[0:0] reshape_simple_add_N_or_3_nl;
  wire[0:0] reshape_simple_add_N_or_15_nl;
  wire[0:0] reshape_simple_add_N_and_3_nl;
  wire[0:0] reshape_simple_add_N_mux1h_5_nl;
  wire[0:0] reshape_simple_add_N_and_4_nl;
  wire[0:0] reshape_simple_add_N_mux1h_6_nl;
  wire[1:0] reshape_simple_add_N_and_5_nl;
  wire[0:0] reshape_simple_add_N_mux1h_7_nl;
  wire[0:0] reshape_simple_add_N_mux1h_10_nl;
  wire[0:0] memory_1_and_nl;
  wire[0:0] memory_1_memory_1_mux_nl;
  wire[13:0] memory_1_and_9_nl;
  wire[13:0] memory_1_mux1h_10_nl;
  wire[13:0] FOR_I_FOR_I_nor_1_nl;
  wire[13:0] BIAS_I_BIAS_I_nor_nl;
  wire[0:0] memory_1_and_10_nl;
  wire[0:0] memory_1_mux1h_11_nl;
  wire[0:0] FOR_I_FOR_I_nor_2_nl;
  wire[0:0] BIAS_I_BIAS_I_nor_3_nl;
  wire[7:0] memory_2_and_3_nl;
  wire[7:0] memory_2_mux1h_1_nl;
  wire[3:0] FOR_B_2_if_acc_12_nl;
  wire[4:0] nl_FOR_B_2_if_acc_12_nl;
  wire[5:0] FOR_B_4_if_acc_16_nl;
  wire[6:0] nl_FOR_B_4_if_acc_16_nl;
  wire[0:0] memory_2_not_4_nl;
  wire[0:0] memory_2_and_4_nl;
  wire[0:0] memory_2_mux1h_4_nl;
  wire[1:0] memory_2_and_5_nl;
  wire[1:0] memory_2_mux1h_5_nl;
  wire[0:0] memory_2_not_6_nl;
  wire[7:0] memory_2_and_nl;
  wire[7:0] memory_2_mux1h_nl;
  wire[3:0] FOR_B_1_if_acc_5_nl;
  wire[4:0] nl_FOR_B_1_if_acc_5_nl;
  wire[5:0] FOR_B_3_if_acc_5_nl;
  wire[6:0] nl_FOR_B_3_if_acc_5_nl;
  wire[0:0] memory_2_not_1_nl;
  wire[0:0] memory_2_and_1_nl;
  wire[0:0] memory_2_mux1h_2_nl;
  wire[1:0] memory_2_and_2_nl;
  wire[1:0] memory_2_mux1h_3_nl;
  wire[0:0] memory_2_not_3_nl;
  wire[15:0] MP1_simple_bigger_mux1h_nl;
  wire[0:0] or_198_nl;
  wire[0:0] memory_2_nand_nl;
  wire[3:0] acc_nl;
  wire[4:0] nl_acc_nl;
  wire[1:0] INIT_I_mux1h_7_nl;
  wire[0:0] INIT_I_or_13_nl;
  wire[0:0] INIT_I_or_14_nl;
  wire[0:0] INIT_I_or_15_nl;
  wire[0:0] INIT_I_nor_1_nl;
  wire[1:0] INIT_I_mux1h_8_nl;
  wire[0:0] INIT_I_or_17_nl;
  wire[3:0] acc_1_nl;
  wire[4:0] nl_acc_1_nl;
  wire[1:0] FOR_A_1_if_mux1h_9_nl;
  wire[2:0] FOR_A_3_if_acc_16_nl;
  wire[3:0] nl_FOR_A_3_if_acc_16_nl;
  wire[0:0] FOR_A_1_if_nor_3_nl;
  wire[0:0] FOR_A_1_if_FOR_A_1_if_or_1_nl;
  wire[1:0] FOR_B_mux1h_6_nl;
  wire[0:0] FOR_B_or_3_nl;
  wire[1:0] FOR_B_FOR_B_mux_1_nl;
  wire[1:0] FOR_B_if_mux1h_6_nl;
  wire[0:0] FOR_B_if_or_4_nl;
  wire[1:0] FOR_B_if_mux1h_7_nl;
  wire[3:0] acc_4_nl;
  wire[4:0] nl_acc_4_nl;
  wire[1:0] FOR_A_1_if_mux1h_10_nl;
  wire[0:0] FOR_A_1_if_and_1_nl;
  wire[1:0] FOR_A_1_if_mux1h_11_nl;
  wire[3:0] FOR_J_1_mux1h_2_nl;
  wire[2:0] FOR_J_3_mux1h_2_nl;
  wire[3:0] FOR_K_6_mux1h_2_nl;
  wire[0:0] FOR_K_6_or_5_nl;
  wire[2:0] mux1h_1_nl;
  wire[0:0] or_nl;
  wire[0:0] or_663_nl;
  wire[0:0] FOR_A_1_if_FOR_A_1_if_and_1_nl;
  wire[1:0] FOR_A_1_if_mux1h_12_nl;
  wire[4:0] INIT_J_mux1h_2_nl;
  wire[4:0] INIT_I_mux1h_9_nl;
  wire[0:0] INIT_I_or_18_nl;
  wire[3:0] INIT_I_mux1h_10_nl;
  wire[3:0] FOR_A_3_if_acc_17_nl;
  wire[4:0] nl_FOR_A_3_if_acc_17_nl;
  wire[0:0] INIT_I_or_19_nl;
  wire[4:0] FOR_B_4_if_mux_2_nl;
  wire[3:0] FOR_B_4_if_mux_3_nl;
  wire[4:0] INIT_I_mux1h_11_nl;
  wire[1:0] INIT_I_mux1h_12_nl;
  wire[5:0] INIT_L_mux1h_2_nl;
  wire[1:0] FOR_B_mux1h_7_nl;
  wire[1:0] FOR_B_mux1h_8_nl;
  wire[4:0] FOR_B_mux1h_9_nl;
  wire[2:0] FOR_B_mux1h_10_nl;
  wire[0:0] FOR_B_or_4_nl;
  wire[1:0] FOR_B_if_mux1h_8_nl;
  wire[0:0] FOR_B_if_mux1h_9_nl;
  wire[31:0] mul_nl;
  wire[15:0] FOR_B_if_mux1h_10_nl;
  wire[15:0] FOR_B_if_mux1h_11_nl;
  wire[0:0] FOR_B_if_or_5_nl;
  wire[3:0] FOR_A_5_if_mux_1_nl;
  wire[17:0] acc_21_nl;
  wire[18:0] nl_acc_21_nl;
  wire[15:0] FOR_I_mux1h_2_nl;
  wire[0:0] FOR_I_or_3_nl;
  wire[0:0] FOR_I_nor_5_nl;
  wire[15:0] FOR_I_mux1h_3_nl;
  wire[0:0] FOR_I_or_5_nl;
  wire[0:0] FOR_B_2_if_mux_4_nl;
  wire[13:0] FOR_B_2_if_mux_5_nl;
  wire[0:0] FOR_B_2_if_mux_6_nl;
  wire[2:0] FOR_A_3_if_mux_2_nl;
  wire[1:0] FOR_A_5_if_acc_21_nl;
  wire[2:0] nl_FOR_A_5_if_acc_21_nl;
  wire[2:0] FOR_A_3_if_mux_3_nl;
  wire[2:0] FOR_B_3_if_mux1h_2_nl;
  wire[1:0] FOR_B_3_if_FOR_B_3_if_mux_1_nl;
  wire[0:0] FOR_B_3_if_or_1_nl;
  wire[2:0] INIT_I_2_mux1h_2_nl;
  wire[1:0] INIT_I_2_mux1h_3_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_INIT_I_C_1_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_INIT_I_C_1_tr0 = ~ reg_INIT_I_slc_INIT_I_acc_2_cse;
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_INIT_J_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_INIT_J_C_0_tr0 = ~ (z_out[2]);
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_INIT_L_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_INIT_L_C_0_tr0 = z_out_13[6];
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_B_C_1_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_B_C_1_tr0 = ~((CR1_simple_b_1_0_sva_1[0])
      ^ (CR1_simple_b_1_0_sva_1[1]));
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_A_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_A_C_0_tr0 = ~((z_out_2[0]) ^ (z_out_2[1]));
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_I_C_2_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_I_C_2_tr0 = ~ FOR_I_slc_FOR_I_acc_2_itm;
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_J_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_J_C_0_tr0 = ~ (z_out[2]);
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_BIAS_I_C_2_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_BIAS_I_C_2_tr0 = ~ BIAS_I_slc_BIAS_I_acc_2_itm;
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_BIAS_J_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_BIAS_J_C_0_tr0 = ~ (z_out[2]);
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_L_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_L_C_0_tr0 = z_out_13[6];
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_A_1_C_1_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_A_1_C_1_tr0 = ~((CR1_simple_b_1_0_sva_1[0])
      ^ (CR1_simple_b_1_0_sva_1[1]));
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_B_1_C_1_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_B_1_C_1_tr0 = ~((CR1_simple_b_1_0_sva_1[0])
      ^ (CR1_simple_b_1_0_sva_1[1]));
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_I_1_C_1_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_I_1_C_1_tr0 = ~ (z_out[2]);
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_J_1_C_1_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_J_1_C_1_tr0 = ~ (z_out[2]);
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_K_1_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_K_1_C_0_tr0 = z_out_13[6];
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_INIT_I_1_C_1_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_INIT_I_1_C_1_tr0 = ~ reg_INIT_I_slc_INIT_I_acc_2_cse;
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_INIT_J_1_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_INIT_J_1_C_0_tr0 = ~ (z_out[2]);
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_INIT_L_1_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_INIT_L_1_C_0_tr0 = z_out_16[5];
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_B_2_C_1_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_B_2_C_1_tr0 = ~((CR1_simple_b_1_0_sva_1[0])
      ^ (CR1_simple_b_1_0_sva_1[1]));
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_A_2_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_A_2_C_0_tr0 = ~((z_out_2[0]) ^
      (z_out_2[1]));
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_I_2_C_2_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_I_2_C_2_tr0 = ~ FOR_I_2_slc_FOR_I_2_acc_2_itm;
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_J_2_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_J_2_C_0_tr0 = ~ (z_out[2]);
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_K_2_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_K_2_C_0_tr0 = z_out_13[6];
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_BIAS_I_1_C_2_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_BIAS_I_1_C_2_tr0 = ~ BIAS_I_1_slc_BIAS_I_1_acc_2_itm;
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_BIAS_J_1_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_BIAS_J_1_C_0_tr0 = ~ (z_out[2]);
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_L_1_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_L_1_C_0_tr0 = z_out_16[5];
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_A_3_C_1_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_A_3_C_1_tr0 = ~((CR1_simple_b_1_0_sva_1[0])
      ^ (CR1_simple_b_1_0_sva_1[1]));
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_B_3_C_1_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_B_3_C_1_tr0 = ~((CR1_simple_b_1_0_sva_1[0])
      ^ (CR1_simple_b_1_0_sva_1[1]));
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_I_3_C_1_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_I_3_C_1_tr0 = ~ (z_out[2]);
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_J_3_C_1_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_J_3_C_1_tr0 = ~ (z_out[2]);
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_K_3_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_K_3_C_0_tr0 = z_out_16[5];
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_INIT_I_2_C_1_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_INIT_I_2_C_1_tr0 = ~ reg_INIT_I_slc_INIT_I_acc_2_cse;
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_INIT_J_2_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_INIT_J_2_C_0_tr0 = ~ (z_out[2]);
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_INIT_L_2_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_INIT_L_2_C_0_tr0 = ~ (z_out_7[3]);
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_B_4_C_1_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_B_4_C_1_tr0 = ~((CR1_simple_b_1_0_sva_1[0])
      ^ (CR1_simple_b_1_0_sva_1[1]));
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_A_4_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_A_4_C_0_tr0 = ~((z_out_2[0]) ^
      (z_out_2[1]));
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_I_4_C_2_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_I_4_C_2_tr0 = ~ FOR_I_4_slc_FOR_I_4_acc_2_itm;
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_J_4_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_J_4_C_0_tr0 = ~ (z_out[2]);
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_K_4_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_K_4_C_0_tr0 = z_out_16[5];
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_BIAS_I_2_C_2_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_BIAS_I_2_C_2_tr0 = ~ BIAS_I_2_slc_BIAS_I_2_acc_2_itm;
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_BIAS_J_2_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_BIAS_J_2_C_0_tr0 = ~ (z_out[2]);
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_L_2_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_L_2_C_0_tr0 = ~ (z_out_7[3]);
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_A_5_C_1_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_A_5_C_1_tr0 = MP3_simple_a_1_0_sva[1];
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_B_5_C_1_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_B_5_C_1_tr0 = ~((CR1_simple_b_1_0_sva_1[0])
      ^ (CR1_simple_b_1_0_sva_1[1]));
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_I_5_C_1_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_I_5_C_1_tr0 = ~((z_out_2[0]) ^
      (z_out_2[1]));
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_J_5_C_1_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_J_5_C_1_tr0 = ~((z_out_2[0]) ^
      (z_out_2[1]));
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_K_5_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_K_5_C_0_tr0 = ~ (z_out_7[3]);
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_K_6_C_2_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_K_6_C_2_tr0 = ~ FOR_K_6_slc_FOR_K_6_acc_3_itm;
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_J_6_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_J_6_C_0_tr0 = ~((z_out_2[0]) ^
      (z_out_2[1]));
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_K_7_C_1_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_K_7_C_1_tr0 = ~ FOR_K_7_slc_FOR_K_7_acc_6_itm;
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_FOR_J_7_C_1_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_FOR_J_7_C_1_tr0 = ~ (z_out_7[3]);
  wire [0:0] nl_CNN_main_simple_core_core_fsm_inst_for_C_0_tr0;
  assign nl_CNN_main_simple_core_core_fsm_inst_for_C_0_tr0 = ~ (z_out_7[3]);
  ccs_out_v1 #(.rscid(32'sd10),
  .width(32'sd4)) index_rsci (
      .idat(index_rsci_idat),
      .dat(index_rsc_dat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) image_rsc_triosy_obj (
      .ld(reg_index_rsc_triosy_obj_ld_cse),
      .lz(image_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) F_1_rsc_triosy_obj (
      .ld(reg_index_rsc_triosy_obj_ld_cse),
      .lz(F_1_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) B_1_rsc_triosy_obj (
      .ld(reg_index_rsc_triosy_obj_ld_cse),
      .lz(B_1_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) F_2_rsc_triosy_obj (
      .ld(reg_index_rsc_triosy_obj_ld_cse),
      .lz(F_2_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) B_2_rsc_triosy_obj (
      .ld(reg_index_rsc_triosy_obj_ld_cse),
      .lz(B_2_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) F_3_rsc_triosy_obj (
      .ld(reg_index_rsc_triosy_obj_ld_cse),
      .lz(F_3_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) B_3_rsc_triosy_obj (
      .ld(reg_index_rsc_triosy_obj_ld_cse),
      .lz(B_3_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) P_W_rsc_triosy_obj (
      .ld(reg_index_rsc_triosy_obj_ld_cse),
      .lz(P_W_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) P_B_rsc_triosy_obj (
      .ld(reg_index_rsc_triosy_obj_ld_cse),
      .lz(P_B_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) index_rsc_triosy_obj (
      .ld(reg_index_rsc_triosy_obj_ld_cse),
      .lz(index_rsc_triosy_lz)
    );
  CNN_main_simple_core_core_fsm CNN_main_simple_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .INIT_I_C_1_tr0(nl_CNN_main_simple_core_core_fsm_inst_INIT_I_C_1_tr0[0:0]),
      .INIT_J_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_INIT_J_C_0_tr0[0:0]),
      .INIT_L_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_INIT_L_C_0_tr0[0:0]),
      .FOR_B_C_1_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_B_C_1_tr0[0:0]),
      .FOR_A_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_A_C_0_tr0[0:0]),
      .FOR_I_C_2_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_I_C_2_tr0[0:0]),
      .FOR_J_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_J_C_0_tr0[0:0]),
      .FOR_K_C_0_tr0(FOR_I_6_FOR_I_6_xnor_cse),
      .BIAS_I_C_2_tr0(nl_CNN_main_simple_core_core_fsm_inst_BIAS_I_C_2_tr0[0:0]),
      .BIAS_J_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_BIAS_J_C_0_tr0[0:0]),
      .FOR_L_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_L_C_0_tr0[0:0]),
      .FOR_A_1_C_1_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_A_1_C_1_tr0[0:0]),
      .FOR_B_1_C_1_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_B_1_C_1_tr0[0:0]),
      .FOR_I_1_C_1_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_I_1_C_1_tr0[0:0]),
      .FOR_J_1_C_1_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_J_1_C_1_tr0[0:0]),
      .FOR_K_1_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_K_1_C_0_tr0[0:0]),
      .INIT_I_1_C_1_tr0(nl_CNN_main_simple_core_core_fsm_inst_INIT_I_1_C_1_tr0[0:0]),
      .INIT_J_1_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_INIT_J_1_C_0_tr0[0:0]),
      .INIT_L_1_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_INIT_L_1_C_0_tr0[0:0]),
      .FOR_B_2_C_1_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_B_2_C_1_tr0[0:0]),
      .FOR_A_2_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_A_2_C_0_tr0[0:0]),
      .FOR_I_2_C_2_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_I_2_C_2_tr0[0:0]),
      .FOR_J_2_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_J_2_C_0_tr0[0:0]),
      .FOR_K_2_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_K_2_C_0_tr0[0:0]),
      .BIAS_I_1_C_2_tr0(nl_CNN_main_simple_core_core_fsm_inst_BIAS_I_1_C_2_tr0[0:0]),
      .BIAS_J_1_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_BIAS_J_1_C_0_tr0[0:0]),
      .FOR_L_1_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_L_1_C_0_tr0[0:0]),
      .FOR_A_3_C_1_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_A_3_C_1_tr0[0:0]),
      .FOR_B_3_C_1_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_B_3_C_1_tr0[0:0]),
      .FOR_I_3_C_1_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_I_3_C_1_tr0[0:0]),
      .FOR_J_3_C_1_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_J_3_C_1_tr0[0:0]),
      .FOR_K_3_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_K_3_C_0_tr0[0:0]),
      .INIT_I_2_C_1_tr0(nl_CNN_main_simple_core_core_fsm_inst_INIT_I_2_C_1_tr0[0:0]),
      .INIT_J_2_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_INIT_J_2_C_0_tr0[0:0]),
      .INIT_L_2_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_INIT_L_2_C_0_tr0[0:0]),
      .FOR_B_4_C_1_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_B_4_C_1_tr0[0:0]),
      .FOR_A_4_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_A_4_C_0_tr0[0:0]),
      .FOR_I_4_C_2_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_I_4_C_2_tr0[0:0]),
      .FOR_J_4_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_J_4_C_0_tr0[0:0]),
      .FOR_K_4_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_K_4_C_0_tr0[0:0]),
      .BIAS_I_2_C_2_tr0(nl_CNN_main_simple_core_core_fsm_inst_BIAS_I_2_C_2_tr0[0:0]),
      .BIAS_J_2_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_BIAS_J_2_C_0_tr0[0:0]),
      .FOR_L_2_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_L_2_C_0_tr0[0:0]),
      .FOR_A_5_C_1_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_A_5_C_1_tr0[0:0]),
      .FOR_B_5_C_1_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_B_5_C_1_tr0[0:0]),
      .FOR_I_5_C_1_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_I_5_C_1_tr0[0:0]),
      .FOR_J_5_C_1_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_J_5_C_1_tr0[0:0]),
      .FOR_K_5_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_K_5_C_0_tr0[0:0]),
      .FOR_K_6_C_2_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_K_6_C_2_tr0[0:0]),
      .FOR_J_6_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_J_6_C_0_tr0[0:0]),
      .FOR_I_6_C_0_tr0(FOR_I_6_FOR_I_6_xnor_cse),
      .FOR_K_7_C_1_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_K_7_C_1_tr0[0:0]),
      .FOR_J_7_C_1_tr0(nl_CNN_main_simple_core_core_fsm_inst_FOR_J_7_C_1_tr0[0:0]),
      .for_C_0_tr0(nl_CNN_main_simple_core_core_fsm_inst_for_C_0_tr0[0:0])
    );
  assign memory_1_or_seb = (fsm_output[68]) | (fsm_output[63]) | (fsm_output[42])
      | (fsm_output[37]) | (fsm_output[16]) | (fsm_output[11]) | (fsm_output[82]);
  assign memory_1_or_1_seb = (fsm_output[68]) | (fsm_output[55]) | (fsm_output[29])
      | (fsm_output[3]) | (fsm_output[63]) | (fsm_output[42]) | (fsm_output[37])
      | (fsm_output[16]) | (fsm_output[11]) | (fsm_output[82]) | (fsm_output[0]);
  assign nand_cse_1 = ~(z_out_1_2 & (z_out[2]));
  assign memory_1_nor_1_seb = ~((~((fsm_output[62]) | (fsm_output[36]) | (fsm_output[10])
      | (fsm_output[67]) | (fsm_output[41]) | (fsm_output[15]) | (fsm_output[74])
      | (fsm_output[48]) | (fsm_output[22]) | (fsm_output[87]))) | (nand_cse_1 &
      (fsm_output[22])) | (nand_cse_1 & (fsm_output[74])) | (nand_cse_1 & (fsm_output[48])));
  assign or_125_cse = FOR_B_oelse_acc_tmp_13 | FOR_B_oelse_2_acc_itm_13;
  assign reg_CR1_simple_l_1_6_0_sva_5_CR1_simple_l_or_cse = (fsm_output[2]) | (fsm_output[6]);
  assign reg_CR1_simple_CR1_simple_aux_or_1_cse = or_332_cse | (fsm_output[9:8]!=2'b00);
  assign or_332_cse = (fsm_output[13]) | (fsm_output[19]) | (fsm_output[14]) | (fsm_output[6])
      | (fsm_output[12]);
  assign reg_CR2_simple_CR2_simple_aux_or_1_cse = or_400_cse | (fsm_output[35:34]!=2'b00);
  assign or_400_cse = (fsm_output[39]) | (fsm_output[45]) | (fsm_output[40]) | (fsm_output[32])
      | (fsm_output[38]);
  assign FOR_B_2_if_FOR_B_2_if_or_cse = FOR_B_2_oelse_2_acc_itm_14 | FOR_B_2_oelse_acc_tmp_14;
  assign reg_CR3_simple_CR3_simple_aux_or_1_cse = or_468_cse | (fsm_output[61:60]!=2'b00);
  assign or_468_cse = (fsm_output[65]) | (fsm_output[71]) | (fsm_output[66]) | (fsm_output[58])
      | (fsm_output[64]);
  assign FOR_B_4_if_FOR_B_4_if_or_cse = (z_out_22[15]) | FOR_B_4_oelse_acc_tmp_15;
  assign reg_MP3_simple_b_1_MP3_simple_b_or_cse = (fsm_output[73]) | (fsm_output[77]);
  assign FOR_J_7_or_29_rgt = (fsm_output[87]) | ((~ FOR_J_7_and_21_cse_sva) & (fsm_output[88]));
  assign FOR_J_7_and_81_rgt = FOR_J_7_and_21_cse_sva & (fsm_output[88]);
  assign FOR_J_7_or_2_rgt = (fsm_output[87]) | ((~ FOR_J_7_and_20_cse_sva) & (fsm_output[88]));
  assign FOR_J_7_and_27_rgt = FOR_J_7_and_20_cse_sva & (fsm_output[88]);
  assign FOR_J_7_or_26_rgt = (fsm_output[87]) | ((~ FOR_J_7_and_19_cse_sva) & (fsm_output[88]));
  assign FOR_J_7_and_75_rgt = FOR_J_7_and_19_cse_sva & (fsm_output[88]);
  assign FOR_J_7_or_23_rgt = (fsm_output[87]) | ((~ FOR_J_7_and_18_cse_sva) & (fsm_output[88]));
  assign FOR_J_7_and_69_rgt = FOR_J_7_and_18_cse_sva & (fsm_output[88]);
  assign FOR_J_7_or_20_rgt = (fsm_output[87]) | ((~ FOR_J_7_and_17_cse_sva) & (fsm_output[88]));
  assign FOR_J_7_and_63_rgt = FOR_J_7_and_17_cse_sva & (fsm_output[88]);
  assign FOR_J_7_or_17_rgt = (fsm_output[87]) | ((~ FOR_J_7_and_16_cse_sva) & (fsm_output[88]));
  assign FOR_J_7_and_57_rgt = FOR_J_7_and_16_cse_sva & (fsm_output[88]);
  assign FOR_J_7_or_14_rgt = (fsm_output[87]) | ((~ FOR_J_7_and_15_cse_sva) & (fsm_output[88]));
  assign FOR_J_7_and_51_rgt = FOR_J_7_and_15_cse_sva & (fsm_output[88]);
  assign FOR_J_7_or_11_rgt = (fsm_output[87]) | ((~ FOR_J_7_and_14_cse_sva) & (fsm_output[88]));
  assign FOR_J_7_and_45_rgt = FOR_J_7_and_14_cse_sva & (fsm_output[88]);
  assign FOR_J_7_or_8_rgt = (fsm_output[87]) | ((~ FOR_J_7_and_13_cse_sva) & (fsm_output[88]));
  assign FOR_J_7_and_39_rgt = FOR_J_7_and_13_cse_sva & (fsm_output[88]);
  assign FOR_J_7_or_5_rgt = (fsm_output[87]) | ((~ FOR_J_7_and_12_cse_sva) & (fsm_output[88]));
  assign FOR_J_7_and_33_rgt = FOR_J_7_and_12_cse_sva & (fsm_output[88]);
  assign CR1_simple_aux_15_lpi_7_mx1 = MUX_s_1_2_2((FOR_B_if_acc_psp_sva_1[18]),
      CR1_simple_aux_15_lpi_7, FOR_B_lor_2_lpi_7_dfm_st);
  assign FOR_B_if_nor_2_nl = ~(MUX_v_14_2_2((FOR_B_if_acc_psp_sva_1[14:1]), 14'b11111111111111,
      FOR_B_if_nor_ovfl_sva_1));
  assign FOR_B_if_FOR_B_if_nor_nl = ~(MUX_v_14_2_2((FOR_B_if_nor_2_nl), 14'b11111111111111,
      FOR_B_if_and_unfl_sva_1));
  assign CR1_simple_aux_14_1_lpi_7_mx1 = MUX_v_14_2_2((FOR_B_if_FOR_B_if_nor_nl),
      CR1_simple_aux_14_1_lpi_7, FOR_B_lor_2_lpi_7_dfm_st);
  assign FOR_B_if_FOR_B_if_nor_1_nl = ~((~((FOR_B_if_acc_psp_sva_1[0]) | FOR_B_if_nor_ovfl_sva_1))
      | FOR_B_if_and_unfl_sva_1);
  assign CR1_simple_aux_0_lpi_7_mx1 = MUX_s_1_2_2((FOR_B_if_FOR_B_if_nor_1_nl), CR1_simple_aux_0_lpi_7,
      FOR_B_lor_2_lpi_7_dfm_st);
  assign nl_FOR_B_if_acc_10_psp_1 = conv_s2u_5_7(FOR_B_if_acc_5_sdt_1[5:1]) + conv_s2u_6_7(FOR_B_acc_1_psp_sva_1);
  assign FOR_B_if_acc_10_psp_1 = nl_FOR_B_if_acc_10_psp_1[6:0];
  assign nl_FOR_B_if_acc_5_sdt_1 = FOR_B_acc_1_psp_sva_1 + conv_s2s_3_6(z_out_16[5:3]);
  assign FOR_B_if_acc_5_sdt_1 = nl_FOR_B_if_acc_5_sdt_1[5:0];
  assign nl_FOR_B_acc_1_psp_sva_1 = conv_s2s_2_6(z_out_15_1_0) + conv_u2s_5_6(CR1_simple_i_2_4_0_sva);
  assign FOR_B_acc_1_psp_sva_1 = nl_FOR_B_acc_1_psp_sva_1[5:0];
  assign nl_FOR_B_oelse_2_acc_nl = ({1'b1 , (signext_13_3(~ (z_out_16[5:3])))}) +
      14'b11;
  assign FOR_B_oelse_2_acc_nl = nl_FOR_B_oelse_2_acc_nl[13:0];
  assign FOR_B_oelse_2_acc_itm_13 = readslicef_14_1_13((FOR_B_oelse_2_acc_nl));
  assign nl_FOR_B_oelse_acc_nl = ({1'b1 , (signext_13_3(~ (FOR_B_acc_1_psp_sva_1[5:3])))})
      + 14'b11;
  assign FOR_B_oelse_acc_nl = nl_FOR_B_oelse_acc_nl[13:0];
  assign FOR_B_oelse_acc_tmp_13 = readslicef_14_1_13((FOR_B_oelse_acc_nl));
  assign nl_FOR_B_if_acc_psp_sva_1 = conv_s2u_16_19({CR1_simple_aux_15_lpi_7 , CR1_simple_aux_14_1_lpi_7
      , CR1_simple_aux_0_lpi_7}) + (z_out_18_31_12[19:1]);
  assign FOR_B_if_acc_psp_sva_1 = nl_FOR_B_if_acc_psp_sva_1[18:0];
  assign FOR_B_if_nor_ovfl_sva_1 = ~((FOR_B_if_acc_psp_sva_1[18]) | (~((FOR_B_if_acc_psp_sva_1[17:15]!=3'b000))));
  assign FOR_B_if_and_unfl_sva_1 = (FOR_B_if_acc_psp_sva_1[18]) & (~((FOR_B_if_acc_psp_sva_1[17:15]==3'b111)));
  assign FOR_I_nor_2_cse = ~((z_out_22[16:15]!=2'b01));
  assign FOR_I_and_4_cse = (z_out_22[16:15]==2'b10);
  assign or_141_cse = reg_FOR_A_1_lor_lpi_6_dfm_cse | (~ (z_out_22[16]));
  assign MP1_simple_bigger_lpi_6_mx1 = MUX_v_16_2_2(memory_1_rsci_q_d, MP1_simple_bigger_lpi_6,
      or_141_cse);
  assign nl_FOR_A_1_oelse_acc_1_ncse_sva_2 = MP1_simple_i_4_1_sva + conv_u2u_1_4(MP1_simple_a_1_0_sva[1]);
  assign FOR_A_1_oelse_acc_1_ncse_sva_2 = nl_FOR_A_1_oelse_acc_1_ncse_sva_2[3:0];
  assign nl_FOR_B_1_if_acc_3_sdt_1 = conv_u2u_6_7(MP1_simple_k_6_0_sva_5_0) + conv_u2u_4_7(z_out_23[4:1]);
  assign FOR_B_1_if_acc_3_sdt_1 = nl_FOR_B_1_if_acc_3_sdt_1[6:0];
  assign CR2_simple_aux_15_lpi_7_mx1 = MUX_s_1_2_2((z_out_24[19]), CR2_simple_aux_15_lpi_7,
      FOR_B_2_lor_2_lpi_7_dfm_st);
  assign FOR_B_2_if_nor_2_nl = ~(MUX_v_14_2_2((z_out_24[14:1]), 14'b11111111111111,
      FOR_B_2_if_nor_ovfl_sva_1));
  assign FOR_B_2_if_FOR_B_2_if_nor_cse = ~(MUX_v_14_2_2((FOR_B_2_if_nor_2_nl), 14'b11111111111111,
      FOR_B_2_if_and_unfl_sva_1));
  assign CR2_simple_aux_14_1_lpi_7_mx1 = MUX_v_14_2_2(FOR_B_2_if_FOR_B_2_if_nor_cse,
      CR2_simple_aux_14_1_lpi_7, FOR_B_2_lor_2_lpi_7_dfm_st);
  assign FOR_B_2_if_FOR_B_2_if_nor_1_cse = ~((~((z_out_24[0]) | FOR_B_2_if_nor_ovfl_sva_1))
      | FOR_B_2_if_and_unfl_sva_1);
  assign CR2_simple_aux_0_lpi_7_mx1 = MUX_s_1_2_2(FOR_B_2_if_FOR_B_2_if_nor_1_cse,
      CR2_simple_aux_0_lpi_7, FOR_B_2_lor_2_lpi_7_dfm_st);
  assign nl_FOR_B_2_if_acc_8_sdt_1 = conv_u2u_6_7(CR2_simple_k_6_0_sva_5_0_1) + conv_s2u_5_7(FOR_B_2_if_acc_9_psp_1[5:1]);
  assign FOR_B_2_if_acc_8_sdt_1 = nl_FOR_B_2_if_acc_8_sdt_1[6:0];
  assign nl_FOR_B_2_if_acc_9_psp_1 = conv_s2u_4_6(z_out_16[4:1]) + conv_s2u_5_6(FOR_B_2_acc_1_psp_sva_1);
  assign FOR_B_2_if_acc_9_psp_1 = nl_FOR_B_2_if_acc_9_psp_1[5:0];
  assign nl_CR2_simple_j_aux_4_0_sva_1 = conv_s2u_2_5(z_out_14_1_0) + conv_u2u_4_5(CR2_simple_j_2_3_0_sva);
  assign CR2_simple_j_aux_4_0_sva_1 = nl_CR2_simple_j_aux_4_0_sva_1[4:0];
  assign nl_FOR_B_2_acc_1_psp_sva_1 = conv_s2s_2_5(z_out_15_1_0) + conv_u2s_4_5(CR2_simple_i_2_3_0_sva);
  assign FOR_B_2_acc_1_psp_sva_1 = nl_FOR_B_2_acc_1_psp_sva_1[4:0];
  assign nl_FOR_B_2_oelse_2_acc_nl = ({1'b1 , (signext_14_3(~ (CR2_simple_j_aux_4_0_sva_1[4:2])))})
      + 15'b11;
  assign FOR_B_2_oelse_2_acc_nl = nl_FOR_B_2_oelse_2_acc_nl[14:0];
  assign FOR_B_2_oelse_2_acc_itm_14 = readslicef_15_1_14((FOR_B_2_oelse_2_acc_nl));
  assign nl_FOR_B_2_oelse_acc_nl = ({1'b1 , (signext_14_3(~ (FOR_B_2_acc_1_psp_sva_1[4:2])))})
      + 15'b11;
  assign FOR_B_2_oelse_acc_nl = nl_FOR_B_2_oelse_acc_nl[14:0];
  assign FOR_B_2_oelse_acc_tmp_14 = readslicef_15_1_14((FOR_B_2_oelse_acc_nl));
  assign FOR_B_2_if_nor_ovfl_sva_1 = ~((z_out_24[19]) | (~((z_out_24[18:15]!=4'b0000))));
  assign FOR_B_2_if_and_unfl_sva_1 = (z_out_24[19]) & (~((z_out_24[18:15]==4'b1111)));
  assign MP2_simple_bigger_lpi_6_mx1 = MUX_v_16_2_2(memory_1_rsci_q_d, MP2_simple_bigger_lpi_6,
      or_141_cse);
  assign nl_FOR_A_3_oelse_acc_1_ncse_sva_2 = MP2_simple_i_3_1_sva + conv_u2u_1_3(MP2_simple_a_1_0_sva[1]);
  assign FOR_A_3_oelse_acc_1_ncse_sva_2 = nl_FOR_A_3_oelse_acc_1_ncse_sva_2[2:0];
  assign nl_FOR_B_3_if_acc_sdt_1 = MP2_simple_j_N_2_0_sva_1 + conv_u2u_2_3(MP2_simple_i_N_2_0_sva_1[2:1]);
  assign FOR_B_3_if_acc_sdt_1 = nl_FOR_B_3_if_acc_sdt_1[2:0];
  assign nl_INIT_I_2_acc_6_sdt_1 = CR3_simple_l_1_4_0_sva + conv_u2u_4_5(z_out_26);
  assign INIT_I_2_acc_6_sdt_1 = nl_INIT_I_2_acc_6_sdt_1[4:0];
  assign CR3_simple_aux_15_lpi_7_mx1 = MUX_s_1_2_2((z_out_24[19]), CR3_simple_aux_15_lpi_7,
      FOR_B_4_lor_2_lpi_7_dfm_st);
  assign CR3_simple_aux_14_1_lpi_7_mx1 = MUX_v_14_2_2(FOR_B_2_if_FOR_B_2_if_nor_cse,
      CR3_simple_aux_14_1_lpi_7, FOR_B_4_lor_2_lpi_7_dfm_st);
  assign CR3_simple_aux_0_lpi_7_mx1 = MUX_s_1_2_2(FOR_B_2_if_FOR_B_2_if_nor_1_cse,
      CR3_simple_aux_0_lpi_7, FOR_B_4_lor_2_lpi_7_dfm_st);
  assign nl_FOR_B_4_if_acc_12_nl = conv_s2s_4_5(FOR_B_4_if_acc_6_sdt_1[4:1]) + conv_s2s_4_5(FOR_B_4_acc_1_psp_1_sva_1);
  assign FOR_B_4_if_acc_12_nl = nl_FOR_B_4_if_acc_12_nl[4:0];
  assign nl_FOR_B_4_if_acc_11_sdt_1 = conv_s2s_5_7(FOR_B_4_if_acc_12_nl) + conv_u2s_5_7(CR3_simple_k_5_0_sva_4_0);
  assign FOR_B_4_if_acc_11_sdt_1 = nl_FOR_B_4_if_acc_11_sdt_1[6:0];
  assign nl_FOR_B_4_if_acc_6_sdt_1 = conv_s2s_4_5(FOR_B_4_acc_1_psp_1_sva_1) + conv_s2s_3_5(CR3_simple_j_aux_3_0_sva_1[3:1]);
  assign FOR_B_4_if_acc_6_sdt_1 = nl_FOR_B_4_if_acc_6_sdt_1[4:0];
  assign nl_CR3_simple_j_aux_3_0_sva_1 = conv_s2u_2_4(z_out_15_1_0) + conv_u2u_3_4(CR3_simple_j_2_2_0_sva);
  assign CR3_simple_j_aux_3_0_sva_1 = nl_CR3_simple_j_aux_3_0_sva_1[3:0];
  assign nl_FOR_B_4_acc_1_psp_1_sva_1 = conv_s2s_2_4(z_out_14_1_0) + conv_u2s_3_4(CR3_simple_i_2_2_0_sva);
  assign FOR_B_4_acc_1_psp_1_sva_1 = nl_FOR_B_4_acc_1_psp_1_sva_1[3:0];
  assign nl_FOR_B_4_if_acc_9_nl = conv_s2s_3_4(z_out) + conv_u2s_3_4(z_out_10[5:3]);
  assign FOR_B_4_if_acc_9_nl = nl_FOR_B_4_if_acc_9_nl[3:0];
  assign nl_FOR_B_4_if_acc_10_sdt_4_0_1 = conv_s2u_4_5(FOR_B_4_if_acc_9_nl) + conv_u2u_4_5({CR3_simple_b_1_0_sva
      , 2'b1});
  assign FOR_B_4_if_acc_10_sdt_4_0_1 = nl_FOR_B_4_if_acc_10_sdt_4_0_1[4:0];
  assign nl_FOR_B_4_oelse_acc_nl = ({1'b1 , (signext_15_3(~ (FOR_B_4_acc_1_psp_1_sva_1[3:1])))})
      + 16'b11;
  assign FOR_B_4_oelse_acc_nl = nl_FOR_B_4_oelse_acc_nl[15:0];
  assign FOR_B_4_oelse_acc_tmp_15 = readslicef_16_1_15((FOR_B_4_oelse_acc_nl));
  assign MP3_simple_bigger_lpi_6_mx1 = MUX_v_16_2_2(memory_1_rsci_q_d, MP3_simple_bigger_lpi_6,
      or_141_cse);
  assign FOR_J_7_and_stg_2_1_sva_1 = FOR_J_7_and_stg_1_1_sva_1 & (~ (perceptron_simple_j_3_0_sva[2]));
  assign FOR_J_7_and_stg_2_0_sva_1 = FOR_J_7_and_stg_1_0_sva_1 & (~ (perceptron_simple_j_3_0_sva[2]));
  assign FOR_J_7_and_stg_1_3_sva_1 = (perceptron_simple_j_3_0_sva[1:0]==2'b11);
  assign FOR_J_7_and_stg_1_2_sva_1 = (perceptron_simple_j_3_0_sva[1:0]==2'b10);
  assign FOR_J_7_and_stg_1_1_sva_1 = (perceptron_simple_j_3_0_sva[1:0]==2'b01);
  assign FOR_J_7_and_stg_1_0_sva_1 = ~((perceptron_simple_j_3_0_sva[1:0]!=2'b00));
  assign nl_perceptron_simple_k_7_0_sva_2 = perceptron_simple_k_7_0_sva + 8'b1;
  assign perceptron_simple_k_7_0_sva_2 = nl_perceptron_simple_k_7_0_sva_2[7:0];
  assign nl_FOR_K_7_acc_8_sdt_1 = perceptron_simple_k_7_0_sva + conv_u2u_3_8(perceptron_simple_j_3_0_sva[3:1]);
  assign FOR_K_7_acc_8_sdt_1 = nl_FOR_K_7_acc_8_sdt_1[7:0];
  assign nl_FOR_K_7_acc_7_psp_sva_1 = conv_s2u_16_17({FOR_K_7_mux_28_itm , FOR_K_7_mux_29_itm
      , FOR_K_7_mux_30_itm}) + (z_out_18_31_12[19:3]);
  assign FOR_K_7_acc_7_psp_sva_1 = nl_FOR_K_7_acc_7_psp_sva_1[16:0];
  assign FOR_K_7_FOR_K_7_nor_2_psp_sva_1 = ~((~((FOR_K_7_acc_7_psp_sva_1[0]) | FOR_K_7_nor_ovfl_sva_1))
      | FOR_K_7_and_unfl_sva_1);
  assign FOR_K_7_nor_3_nl = ~(MUX_v_14_2_2((FOR_K_7_acc_7_psp_sva_1[14:1]), 14'b11111111111111,
      FOR_K_7_nor_ovfl_sva_1));
  assign FOR_K_7_FOR_K_7_nor_1_psp_sva_1 = ~(MUX_v_14_2_2((FOR_K_7_nor_3_nl), 14'b11111111111111,
      FOR_K_7_and_unfl_sva_1));
  assign FOR_K_7_nor_ovfl_sva_1 = ~((FOR_K_7_acc_7_psp_sva_1[16:15]!=2'b01));
  assign FOR_K_7_and_unfl_sva_1 = (FOR_K_7_acc_7_psp_sva_1[16:15]==2'b10);
  assign max_sva_14_1_mx1 = MUX_v_14_2_2(max_sva_14_1, for_slc_Prob_16_15_0_cse_sva_14_1_1,
      z_out_22[16]);
  assign for_slc_Prob_16_15_0_cse_sva_14_1_1 = MUX_v_14_10_2(Prob_0_sva_2_14_1, Prob_1_14_1_sva_2,
      Prob_2_14_1_sva_2, Prob_3_14_1_sva_2, Prob_4_14_1_sva_2, Prob_5_14_1_sva_2,
      Prob_6_14_1_sva_2, Prob_7_14_1_sva_2, Prob_8_14_1_sva_2, Prob_9_14_1_sva_2,
      k_sva);
  assign for_slc_Prob_16_15_0_cse_sva_15_1 = MUX_s_1_10_2(Prob_0_sva_2_15, Prob_1_15_sva_2,
      Prob_2_15_sva_2, Prob_3_15_sva_2, Prob_4_15_sva_2, Prob_5_15_sva_2, Prob_6_15_sva_2,
      Prob_7_15_sva_2, Prob_8_15_sva_2, Prob_9_15_sva_2, k_sva);
  assign for_slc_Prob_16_15_0_cse_sva_0_1 = MUX_s_1_10_2(Prob_0_sva_2_0, Prob_1_0_sva_2,
      Prob_2_0_sva_2, Prob_3_0_sva_2, Prob_4_0_sva_2, Prob_5_0_sva_2, Prob_6_0_sva_2,
      Prob_7_0_sva_2, Prob_8_0_sva_2, Prob_9_0_sva_2, k_sva);
  assign FOR_I_6_FOR_I_6_xnor_cse = ~((z_out_2[0]) ^ (z_out_2[1]));
  assign and_4_cse = (fsm_output[10:9]!=2'b00);
  assign and_10_cse = (fsm_output[36:35]!=2'b00);
  assign and_16_cse = (fsm_output[62:61]!=2'b00);
  assign or_dcpl_53 = (fsm_output[1]) | (fsm_output[91]);
  assign and_dcpl_6 = ~((fsm_output[76]) | (fsm_output[50]));
  assign and_dcpl_133 = (perceptron_simple_j_3_0_sva[3:2]==2'b10);
  assign or_dcpl_130 = (perceptron_simple_j_3_0_sva[1:0]!=2'b01);
  assign or_dcpl_131 = (perceptron_simple_j_3_0_sva[3:2]!=2'b10);
  assign and_dcpl_136 = ~((perceptron_simple_j_3_0_sva[3:2]!=2'b00));
  assign or_dcpl_134 = (perceptron_simple_j_3_0_sva[1:0]!=2'b00);
  assign or_dcpl_135 = (perceptron_simple_j_3_0_sva[3:2]!=2'b00);
  assign and_dcpl_141 = (perceptron_simple_j_3_0_sva[3:2]==2'b01);
  assign or_dcpl_139 = ~((perceptron_simple_j_3_0_sva[1:0]==2'b11));
  assign or_dcpl_140 = (perceptron_simple_j_3_0_sva[3:2]!=2'b01);
  assign or_dcpl_142 = (perceptron_simple_j_3_0_sva[1:0]!=2'b10);
  assign and_285_cse = (~(FOR_B_2_oelse_acc_tmp_14 | FOR_B_2_oelse_2_acc_itm_14))
      & (fsm_output[33]);
  assign and_283_cse = (~(FOR_B_4_oelse_acc_tmp_15 | (z_out_22[15]))) & (fsm_output[59]);
  assign and_307_cse = FOR_B_2_if_FOR_B_2_if_or_cse & (fsm_output[33]);
  assign and_316_cse = z_out_1_2 & (z_out[2]) & (fsm_output[22]);
  assign and_318_cse = z_out_1_2 & (z_out[2]) & (fsm_output[48]);
  assign and_317_cse = z_out_1_2 & (z_out[2]) & (fsm_output[74]);
  assign and_386_cse = (z_out_7[3]) & (fsm_output[89]);
  assign or_tmp_111 = (~((fsm_output[33]) | (fsm_output[0]))) | and_307_cse;
  assign or_tmp_117 = (~(FOR_B_oelse_acc_tmp_13 | FOR_B_oelse_2_acc_itm_13)) & (fsm_output[7]);
  assign or_tmp_125 = ~((fsm_output[88:86]!=3'b000));
  assign or_tmp_376 = (fsm_output[90:89]!=2'b00);
  assign or_tmp_379 = and_dcpl_133 & FOR_J_7_and_stg_1_1_sva_1 & (fsm_output[86]);
  assign or_tmp_380 = (or_dcpl_131 | or_dcpl_130) & (fsm_output[86]);
  assign or_tmp_383 = (fsm_output[88:87]!=2'b00);
  assign or_tmp_392 = and_dcpl_136 & FOR_J_7_and_stg_1_0_sva_1 & (fsm_output[86]);
  assign or_tmp_393 = (or_dcpl_135 | or_dcpl_134) & (fsm_output[86]);
  assign or_tmp_405 = and_dcpl_133 & FOR_J_7_and_stg_1_0_sva_1 & (fsm_output[86]);
  assign or_tmp_406 = (or_dcpl_131 | or_dcpl_134) & (fsm_output[86]);
  assign or_tmp_418 = and_dcpl_136 & FOR_J_7_and_stg_1_1_sva_1 & (fsm_output[86]);
  assign or_tmp_419 = (or_dcpl_135 | or_dcpl_130) & (fsm_output[86]);
  assign or_tmp_431 = and_dcpl_141 & FOR_J_7_and_stg_1_3_sva_1 & (fsm_output[86]);
  assign or_tmp_432 = (or_dcpl_140 | or_dcpl_139) & (fsm_output[86]);
  assign or_tmp_444 = and_dcpl_136 & FOR_J_7_and_stg_1_2_sva_1 & (fsm_output[86]);
  assign or_tmp_445 = (or_dcpl_135 | or_dcpl_142) & (fsm_output[86]);
  assign or_tmp_457 = and_dcpl_141 & FOR_J_7_and_stg_1_2_sva_1 & (fsm_output[86]);
  assign or_tmp_458 = (or_dcpl_140 | or_dcpl_142) & (fsm_output[86]);
  assign or_tmp_470 = and_dcpl_136 & FOR_J_7_and_stg_1_3_sva_1 & (fsm_output[86]);
  assign or_tmp_471 = (or_dcpl_135 | or_dcpl_139) & (fsm_output[86]);
  assign or_tmp_483 = and_dcpl_141 & FOR_J_7_and_stg_1_1_sva_1 & (fsm_output[86]);
  assign or_tmp_484 = (or_dcpl_140 | or_dcpl_130) & (fsm_output[86]);
  assign or_tmp_496 = and_dcpl_141 & FOR_J_7_and_stg_1_0_sva_1 & (fsm_output[86]);
  assign or_tmp_497 = (or_dcpl_140 | or_dcpl_134) & (fsm_output[86]);
  assign memory_2_rsci_wadr_d_mx0c0 = and_dcpl_6 & (~ (fsm_output[24]));
  assign memory_2_rsci_radr_d_mx0c0 = (~((fsm_output[81]) | (fsm_output[59]) | (fsm_output[33])))
      | (FOR_B_4_if_FOR_B_4_if_or_cse & (fsm_output[59])) | and_307_cse;
  assign reshape_simple_add_N_10_0_lpi_4_mx0c1 = (fsm_output[85:83]!=3'b000);
  assign nl_INIT_I_asn_CR1_simple_add_AF_10_INIT_I_acc_sdt = ({z_out_17 , (z_out_10[4:2])})
      + (CR1_simple_l_1_6_0_sva_5_0[4:0]);
  assign INIT_I_asn_CR1_simple_add_AF_10_INIT_I_acc_sdt = nl_INIT_I_asn_CR1_simple_add_AF_10_INIT_I_acc_sdt[4:0];
  assign or_220_ssc = (fsm_output[82]) | (fsm_output[0]);
  assign nl_FOR_A_1_if_asn_MP1_simple_add_M_10_FOR_A_1_if_acc_sdt = ({z_out_17 ,
      (z_out_23[3:1])}) + (MP1_simple_k_6_0_sva_5_0[4:0]);
  assign FOR_A_1_if_asn_MP1_simple_add_M_10_FOR_A_1_if_acc_sdt = nl_FOR_A_1_if_asn_MP1_simple_add_M_10_FOR_A_1_if_acc_sdt[4:0];
  assign nl_FOR_B_if_asn_CR1_simple_add_M_10_FOR_B_if_acc_nl = ({CR1_simple_k_1_0_sva
      , 1'b0 , CR1_simple_k_1_0_sva}) + (FOR_B_if_acc_10_psp_1[6:2]);
  assign FOR_B_if_asn_CR1_simple_add_M_10_FOR_B_if_acc_nl = nl_FOR_B_if_asn_CR1_simple_add_M_10_FOR_B_if_acc_nl[4:0];
  assign BIAS_I_BIAS_I_and_2_nl = MUX_v_5_2_2(5'b00000, (FOR_B_if_asn_CR1_simple_add_M_10_FOR_B_if_acc_nl),
      or_tmp_117);
  assign FOR_K_FOR_K_and_5_nl = MUX_v_2_2_2(2'b00, (FOR_B_if_acc_10_psp_1[1:0]),
      or_tmp_117);
  assign BIAS_I_BIAS_I_and_3_nl = (FOR_B_if_acc_5_sdt_1[0]) & or_tmp_117;
  assign BIAS_I_2_BIAS_I_2_and_3_nl = MUX_v_3_2_2(3'b000, (z_out_16[2:0]), or_tmp_117);
  assign image_rsci_radr_d = {(BIAS_I_BIAS_I_and_2_nl) , (FOR_K_FOR_K_and_5_nl) ,
      (BIAS_I_BIAS_I_and_3_nl) , (BIAS_I_2_BIAS_I_2_and_3_nl)};
  assign image_rsci_re_d_pff = or_tmp_117;
  assign FOR_K_FOR_K_and_4_nl = (((z_out_7[3]) & (CR1_simple_a_1_0_sva[0])) ^ (CR1_simple_a_1_0_sva[1]))
      & or_tmp_117;
  assign FOR_K_FOR_K_and_11_nl = ((z_out_7[3]) ^ (CR1_simple_a_1_0_sva[0])) & or_tmp_117;
  assign BIAS_I_2_BIAS_I_2_and_2_nl = MUX_v_3_2_2(3'b000, (z_out_7[2:0]), or_tmp_117);
  assign CR1_simple_l_nor_nl = ~((~((fsm_output[7]) | (fsm_output[0]))) | (or_125_cse
      & (fsm_output[7])));
  assign CR1_simple_l_CR1_simple_l_and_1_nl = MUX_v_6_2_2(6'b000000, CR1_simple_l_6_0_sva_5_0_1,
      (CR1_simple_l_nor_nl));
  assign F_1_rsci_radr_d = {(FOR_K_FOR_K_and_4_nl) , (FOR_K_FOR_K_and_11_nl) , (BIAS_I_2_BIAS_I_2_and_2_nl)
      , (CR1_simple_l_CR1_simple_l_and_1_nl)};
  assign B_1_nor_nl = ~((~((fsm_output[17]) | (fsm_output[18]) | (fsm_output[14])
      | (fsm_output[0]))) | ((~ BIAS_I_slc_BIAS_I_acc_2_itm) & (fsm_output[17]))
      | (((z_out_2[0]) ^ (z_out_2[1])) & (fsm_output[14])) | ((~ (z_out[2])) & (fsm_output[18])));
  assign B_1_rsci_radr_d = MUX_v_6_2_2(6'b000000, CR1_simple_l_6_0_sva_5_0_1, (B_1_nor_nl));
  assign B_1_rsci_re_d = (BIAS_I_slc_BIAS_I_acc_2_itm & (fsm_output[17])) | (FOR_I_6_FOR_I_6_xnor_cse
      & (fsm_output[14])) | ((z_out[2]) & (fsm_output[18]));
  assign BIAS_I_2_BIAS_I_2_and_1_nl = MUX_v_3_2_2(3'b000, z_out_3, and_285_cse);
  assign BIAS_I_BIAS_I_and_1_nl = (z_out_4[0]) & and_285_cse;
  assign CR2_simple_k_not_nl = ~ or_tmp_111;
  assign CR2_simple_k_CR2_simple_k_and_nl = MUX_v_6_2_2(6'b000000, CR2_simple_k_6_0_sva_5_0_1,
      (CR2_simple_k_not_nl));
  assign CR2_simple_l_not_nl = ~ or_tmp_111;
  assign CR2_simple_l_CR2_simple_l_and_1_nl = MUX_v_5_2_2(5'b00000, CR2_simple_l_5_0_sva_4_0_1,
      (CR2_simple_l_not_nl));
  assign F_2_rsci_radr_d = {(BIAS_I_2_BIAS_I_2_and_1_nl) , (BIAS_I_BIAS_I_and_1_nl)
      , (CR2_simple_k_CR2_simple_k_and_nl) , (CR2_simple_l_CR2_simple_l_and_1_nl)};
  assign F_2_rsci_re_d = and_285_cse;
  assign B_2_nor_nl = ~((~((fsm_output[43]) | (fsm_output[44]) | (fsm_output[40])
      | (fsm_output[0]))) | ((~ BIAS_I_1_slc_BIAS_I_1_acc_2_itm) & (fsm_output[43]))
      | ((~ (z_out[2])) & (fsm_output[44])) | ((~ (z_out_13[6])) & (fsm_output[40])));
  assign B_2_rsci_radr_d = MUX_v_5_2_2(5'b00000, CR2_simple_l_5_0_sva_4_0_1, (B_2_nor_nl));
  assign B_2_rsci_re_d = (BIAS_I_1_slc_BIAS_I_1_acc_2_itm & (fsm_output[43])) | ((z_out[2])
      & (fsm_output[44])) | ((z_out_13[6]) & (fsm_output[40]));
  assign FOR_K_FOR_K_and_3_nl = (((FOR_B_4_if_acc_10_sdt_4_0_1[4]) & (CR3_simple_a_1_0_sva[0]))
      ^ (FOR_B_4_if_acc_10_sdt_4_0_1[4]) ^ (CR3_simple_a_1_0_sva[1])) & and_283_cse;
  assign FOR_K_FOR_K_and_10_nl = ((FOR_B_4_if_acc_10_sdt_4_0_1[4]) ^ (CR3_simple_a_1_0_sva[0]))
      & and_283_cse;
  assign BIAS_I_1_BIAS_I_1_and_nl = MUX_v_4_2_2(4'b0000, (FOR_B_4_if_acc_10_sdt_4_0_1[3:0]),
      and_283_cse);
  assign BIAS_I_2_BIAS_I_2_and_nl = MUX_v_3_2_2(3'b000, (z_out_10[2:0]), and_283_cse);
  assign FOR_K_FOR_K_and_2_nl = MUX_v_2_2_2(2'b00, (z_out_11[1:0]), and_283_cse);
  assign FOR_K_FOR_K_and_1_nl = MUX_v_2_2_2(2'b00, (CR3_simple_l_4_0_sva[1:0]), and_283_cse);
  assign F_3_rsci_radr_d = {(FOR_K_FOR_K_and_3_nl) , (FOR_K_FOR_K_and_10_nl) , (BIAS_I_1_BIAS_I_1_and_nl)
      , (BIAS_I_2_BIAS_I_2_and_nl) , (FOR_K_FOR_K_and_2_nl) , (FOR_K_FOR_K_and_1_nl)};
  assign F_3_rsci_re_d = and_283_cse;
  assign B_3_nor_nl = ~((~((fsm_output[69]) | (fsm_output[70]) | (fsm_output[66])
      | (fsm_output[0]))) | ((~ BIAS_I_2_slc_BIAS_I_2_acc_2_itm) & (fsm_output[69]))
      | ((~ (z_out[2])) & (fsm_output[70])) | ((~ (z_out_16[5])) & (fsm_output[66])));
  assign B_3_rsci_radr_d = MUX_v_5_2_2(5'b00000, CR3_simple_l_4_0_sva, (B_3_nor_nl));
  assign B_3_rsci_re_d = (BIAS_I_2_slc_BIAS_I_2_acc_2_itm & (fsm_output[69])) | ((z_out[2])
      & (fsm_output[70])) | ((z_out_16[5]) & (fsm_output[66]));
  assign nl_FOR_K_7_acc_9_nl = conv_u2u_6_8(FOR_K_7_acc_8_sdt_1[7:2]) + perceptron_simple_k_7_0_sva;
  assign FOR_K_7_acc_9_nl = nl_FOR_K_7_acc_9_nl[7:0];
  assign FOR_K_7_FOR_K_7_and_nl = MUX_v_8_2_2(8'b00000000, (FOR_K_7_acc_9_nl), (fsm_output[87]));
  assign FOR_K_FOR_K_and_nl = MUX_v_2_2_2(2'b00, (FOR_K_7_acc_8_sdt_1[1:0]), (fsm_output[87]));
  assign BIAS_I_BIAS_I_and_nl = (perceptron_simple_j_3_0_sva[0]) & (fsm_output[87]);
  assign P_W_rsci_radr_d = {(FOR_K_7_FOR_K_7_and_nl) , (FOR_K_FOR_K_and_nl) , (BIAS_I_BIAS_I_and_nl)};
  assign P_W_rsci_re_d = fsm_output[87];
  assign P_B_rsci_radr_d = MUX_v_4_2_2(4'b0000, z_out_5, and_386_cse);
  assign P_B_rsci_re_d = (FOR_I_6_FOR_I_6_xnor_cse & (fsm_output[85])) | and_386_cse;
  assign memory_1_or_2_cse = (fsm_output[10]) | (fsm_output[15]);
  assign memory_1_or_5_cse = (fsm_output[36]) | (fsm_output[41]);
  assign memory_1_or_6_cse_1 = (fsm_output[62]) | (fsm_output[67]);
  assign memory_1_or_3_cse = (fsm_output[36]) | (fsm_output[41]) | and_318_cse;
  assign memory_1_or_12_cse = (fsm_output[62]) | (fsm_output[67]) | and_317_cse;
  assign memory_1_or_13_cse = (fsm_output[10]) | (fsm_output[15]) | (fsm_output[36])
      | (fsm_output[41]) | and_318_cse;
  assign memory_1_mux1h_1_nl = MUX1HOT_s_1_3_2((z_out_19[4]), (FOR_A_1_if_asn_MP1_simple_add_M_10_FOR_A_1_if_acc_sdt[4]),
      (z_out_7[3]), {memory_1_or_2_cse , and_316_cse , memory_1_or_3_cse});
  assign memory_1_and_1_nl = (memory_1_mux1h_1_nl) & (~((fsm_output[62]) | (fsm_output[67])
      | and_317_cse | (fsm_output[87]))) & memory_1_nor_1_seb;
  assign memory_1_mux1h_5_nl = MUX1HOT_v_4_5_2((z_out_19[3:0]), (FOR_A_1_if_asn_MP1_simple_add_M_10_FOR_A_1_if_acc_sdt[3:0]),
      ({(z_out_7[2:0]) , (z_out_10[2])}), (z_out_12[4:1]), ({2'b0 , (perceptron_simple_k_7_0_sva[7:6])}),
      {memory_1_or_2_cse , and_316_cse , memory_1_or_3_cse , memory_1_or_12_cse ,
      (fsm_output[87])});
  assign memory_1_mux1h_12_nl = MUX1HOT_s_1_4_2((z_out_10[1]), (z_out_23[0]), (z_out_12[0]),
      (perceptron_simple_k_7_0_sva[5]), {memory_1_or_13_cse , and_316_cse , memory_1_or_12_cse
      , (fsm_output[87])});
  assign memory_1_mux1h_13_nl = MUX1HOT_s_1_5_2((z_out_10[0]), (z_out_8[0]), (z_out_20[2]),
      (z_out_21[2]), (perceptron_simple_k_7_0_sva[4]), {memory_1_or_13_cse , and_316_cse
      , memory_1_or_6_cse_1 , and_317_cse , (fsm_output[87])});
  assign memory_1_and_4_nl = MUX_v_6_2_2(6'b000000, ({(memory_1_mux1h_5_nl) , (memory_1_mux1h_12_nl)
      , (memory_1_mux1h_13_nl)}), memory_1_nor_1_seb);
  assign memory_1_mux1h_6_nl = MUX1HOT_s_1_7_2((z_out_12[0]), (z_out_4[0]), (z_out_23[0]),
      (z_out_25[0]), (z_out_20[1]), (z_out_21[1]), (perceptron_simple_k_7_0_sva[3]),
      {memory_1_or_2_cse , and_316_cse , memory_1_or_5_cse , and_318_cse , memory_1_or_6_cse_1
      , and_317_cse , (fsm_output[87])});
  assign memory_1_and_5_nl = (memory_1_mux1h_6_nl) & memory_1_nor_1_seb;
  assign memory_1_mux1h_7_nl = MUX1HOT_s_1_8_2((CR1_simple_j_2_4_0_sva[2]), (CR1_simple_j_4_0_sva[2]),
      (FOR_A_1_oelse_acc_1_ncse_sva_2[1]), (z_out_8[0]), (z_out_4[0]), (z_out_20[0]),
      (z_out_21[0]), (perceptron_simple_k_7_0_sva[2]), {(fsm_output[10]) , (fsm_output[15])
      , and_316_cse , memory_1_or_5_cse , and_318_cse , memory_1_or_6_cse_1 , and_317_cse
      , (fsm_output[87])});
  assign memory_1_and_6_nl = (memory_1_mux1h_7_nl) & memory_1_nor_1_seb;
  assign memory_1_mux1h_8_nl = MUX1HOT_s_1_9_2((CR1_simple_j_2_4_0_sva[1]), (CR1_simple_j_4_0_sva[1]),
      (FOR_A_1_oelse_acc_1_ncse_sva_2[0]), (CR2_simple_j_2_3_0_sva[1]), (CR2_simple_j_3_0_sva[1]),
      (FOR_A_3_oelse_acc_1_ncse_sva_2[0]), (z_out_27_2_0[0]), (z_out_4[0]), (perceptron_simple_k_7_0_sva[1]),
      {(fsm_output[10]) , (fsm_output[15]) , and_316_cse , (fsm_output[36]) , (fsm_output[41])
      , and_318_cse , memory_1_or_6_cse_1 , and_317_cse , (fsm_output[87])});
  assign memory_1_and_7_nl = (memory_1_mux1h_8_nl) & memory_1_nor_1_seb;
  assign memory_1_mux1h_9_nl = MUX1HOT_s_1_10_2((CR1_simple_j_2_4_0_sva[0]), (CR1_simple_j_4_0_sva[0]),
      (MP1_simple_a_1_0_sva[0]), (CR2_simple_j_2_3_0_sva[0]), (CR2_simple_j_3_0_sva[0]),
      (MP2_simple_a_1_0_sva[0]), (CR3_simple_j_2_2_0_sva[0]), (CR3_simple_j_2_0_sva[0]),
      (MP3_simple_a_1_0_sva[0]), (perceptron_simple_k_7_0_sva[0]), {(fsm_output[10])
      , (fsm_output[15]) , and_316_cse , (fsm_output[36]) , (fsm_output[41]) , and_318_cse
      , (fsm_output[62]) , (fsm_output[67]) , and_317_cse , (fsm_output[87])});
  assign memory_1_and_8_nl = (memory_1_mux1h_9_nl) & memory_1_nor_1_seb;
  assign memory_1_rsci_radr_d = {(memory_1_and_1_nl) , (memory_1_and_4_nl) , (memory_1_and_5_nl)
      , (memory_1_and_6_nl) , (memory_1_and_7_nl) , (memory_1_and_8_nl)};
  assign reshape_simple_add_N_or_cse = (fsm_output[11]) | (fsm_output[16]);
  assign reshape_simple_add_N_or_11_cse = (fsm_output[37]) | (fsm_output[42]);
  assign reshape_simple_add_N_or_2_cse = (fsm_output[63]) | (fsm_output[68]);
  assign reshape_simple_add_N_mux1h_nl = MUX1HOT_s_1_5_2((reshape_simple_add_N_10_0_lpi_4[10]),
      (INIT_I_asn_CR1_simple_add_AF_10_INIT_I_acc_sdt[4]), (reg_FOR_I_asn_CR1_simple_add_AF_10_FOR_I_acc_psp_cse[4]),
      (z_out_7[3]), (reg_FOR_I_2_acc_11_psp_cse[3]), {or_220_ssc , (fsm_output[3])
      , reshape_simple_add_N_or_cse , (fsm_output[29]) , reshape_simple_add_N_or_11_cse});
  assign reshape_simple_add_N_and_nl = (reshape_simple_add_N_mux1h_nl) & (~((fsm_output[55])
      | (fsm_output[63]) | (fsm_output[68]))) & memory_1_or_1_seb;
  assign reshape_simple_add_N_mux1h_4_nl = MUX1HOT_v_4_7_2((reshape_simple_add_N_10_0_lpi_4[9:6]),
      (INIT_I_asn_CR1_simple_add_AF_10_INIT_I_acc_sdt[3:0]), (reg_FOR_I_asn_CR1_simple_add_AF_10_FOR_I_acc_psp_cse[3:0]),
      ({(z_out_7[2:0]) , (z_out_10[2])}), ({(reg_FOR_I_2_acc_11_psp_cse[2:0]) , (reg_FOR_I_2_acc_9_sdt_cse[2])}),
      (z_out_12[4:1]), (reg_FOR_I_4_acc_11_psp_cse[4:1]), {or_220_ssc , (fsm_output[3])
      , reshape_simple_add_N_or_cse , (fsm_output[29]) , reshape_simple_add_N_or_11_cse
      , (fsm_output[55]) , reshape_simple_add_N_or_2_cse});
  assign reshape_simple_add_N_or_3_nl = (fsm_output[3]) | (fsm_output[29]);
  assign reshape_simple_add_N_or_15_nl = reshape_simple_add_N_or_cse | reshape_simple_add_N_or_11_cse;
  assign reshape_simple_add_N_mux1h_9_nl = MUX1HOT_v_2_5_2((reshape_simple_add_N_10_0_lpi_4[5:4]),
      (z_out_10[1:0]), (reg_FOR_I_2_acc_9_sdt_cse[1:0]), ({(z_out_12[0]) , (INIT_I_2_acc_6_sdt_1[2])}),
      ({(reg_FOR_I_4_acc_11_psp_cse[0]) , (reg_FOR_I_4_acc_9_sdt_cse[2])}), {or_220_ssc
      , (reshape_simple_add_N_or_3_nl) , (reshape_simple_add_N_or_15_nl) , (fsm_output[55])
      , reshape_simple_add_N_or_2_cse});
  assign reshape_simple_add_N_and_2_nl = MUX_v_6_2_2(6'b000000, ({(reshape_simple_add_N_mux1h_4_nl)
      , (reshape_simple_add_N_mux1h_9_nl)}), memory_1_or_1_seb);
  assign reshape_simple_add_N_mux1h_5_nl = MUX1HOT_s_1_7_2((reshape_simple_add_N_10_0_lpi_4[3]),
      (z_out_12[0]), (reg_FOR_I_4_acc_11_psp_cse[0]), (z_out_23[0]), reg_FOR_I_2_acc_10_psp_cse,
      (INIT_I_2_acc_6_sdt_1[1]), (reg_FOR_I_4_acc_9_sdt_cse[1]), {or_220_ssc , (fsm_output[3])
      , reshape_simple_add_N_or_cse , (fsm_output[29]) , reshape_simple_add_N_or_11_cse
      , (fsm_output[55]) , reshape_simple_add_N_or_2_cse});
  assign reshape_simple_add_N_and_3_nl = (reshape_simple_add_N_mux1h_5_nl) & memory_1_or_1_seb;
  assign reshape_simple_add_N_mux1h_6_nl = MUX1HOT_s_1_8_2((reshape_simple_add_N_10_0_lpi_4[2]),
      (CR1_simple_j_1_4_0_sva[2]), (CR1_simple_j_2_4_0_sva[2]), (CR1_simple_j_4_0_sva[2]),
      (z_out_8[0]), reg_FOR_I_2_acc_8_sdt_cse, (INIT_I_2_acc_6_sdt_1[0]), (reg_FOR_I_4_acc_9_sdt_cse[0]),
      {or_220_ssc , (fsm_output[3]) , (fsm_output[11]) , (fsm_output[16]) , (fsm_output[29])
      , reshape_simple_add_N_or_11_cse , (fsm_output[55]) , reshape_simple_add_N_or_2_cse});
  assign reshape_simple_add_N_and_4_nl = (reshape_simple_add_N_mux1h_6_nl) & memory_1_or_1_seb;
  assign reshape_simple_add_N_mux1h_7_nl = MUX1HOT_s_1_9_2((reshape_simple_add_N_10_0_lpi_4[1]),
      (CR1_simple_j_1_4_0_sva[1]), (CR1_simple_j_2_4_0_sva[1]), (CR1_simple_j_4_0_sva[1]),
      (CR2_simple_j_1_3_0_sva[1]), (CR2_simple_j_2_3_0_sva[1]), (CR2_simple_j_3_0_sva[1]),
      (z_out_27_2_0[0]), reg_FOR_I_4_acc_8_sdt_2_0_cse, {or_220_ssc , (fsm_output[3])
      , (fsm_output[11]) , (fsm_output[16]) , (fsm_output[29]) , (fsm_output[37])
      , (fsm_output[42]) , (fsm_output[55]) , reshape_simple_add_N_or_2_cse});
  assign reshape_simple_add_N_mux1h_10_nl = MUX1HOT_s_1_10_2((reshape_simple_add_N_10_0_lpi_4[0]),
      (CR1_simple_j_1_4_0_sva[0]), (CR1_simple_j_2_4_0_sva[0]), (CR1_simple_j_4_0_sva[0]),
      (CR2_simple_j_1_3_0_sva[0]), (CR2_simple_j_2_3_0_sva[0]), (CR2_simple_j_3_0_sva[0]),
      (CR3_simple_j_1_2_0_sva[0]), (CR3_simple_j_2_2_0_sva[0]), (CR3_simple_j_2_0_sva[0]),
      {or_220_ssc , (fsm_output[3]) , (fsm_output[11]) , (fsm_output[16]) , (fsm_output[29])
      , (fsm_output[37]) , (fsm_output[42]) , (fsm_output[55]) , (fsm_output[63])
      , (fsm_output[68])});
  assign reshape_simple_add_N_and_5_nl = MUX_v_2_2_2(2'b00, ({(reshape_simple_add_N_mux1h_7_nl)
      , (reshape_simple_add_N_mux1h_10_nl)}), memory_1_or_1_seb);
  assign memory_1_rsci_wadr_d = {(reshape_simple_add_N_and_nl) , (reshape_simple_add_N_and_2_nl)
      , (reshape_simple_add_N_and_3_nl) , (reshape_simple_add_N_and_4_nl) , (reshape_simple_add_N_and_5_nl)};
  assign FOR_I_nor_3_cse = ~(MUX_v_14_2_2((z_out_22[14:1]), 14'b11111111111111, FOR_I_nor_2_cse));
  assign FOR_I_nor_4_cse = ~((z_out_22[0]) | FOR_I_nor_2_cse);
  assign memory_1_or_17_cse = (fsm_output[11]) | (fsm_output[37]) | (fsm_output[63]);
  assign memory_1_or_19_cse = (fsm_output[16]) | (fsm_output[42]) | (fsm_output[68]);
  assign memory_1_memory_1_mux_nl = MUX_s_1_2_2((z_out_22[16]), (memory_2_rsci_q_d[15]),
      fsm_output[82]);
  assign memory_1_and_nl = (memory_1_memory_1_mux_nl) & (~((fsm_output[16]) | (fsm_output[42])
      | (fsm_output[68]))) & memory_1_or_seb;
  assign FOR_I_FOR_I_nor_1_nl = ~(MUX_v_14_2_2(FOR_I_nor_3_cse, 14'b11111111111111,
      FOR_I_and_4_cse));
  assign BIAS_I_BIAS_I_nor_nl = ~(FOR_I_nor_3_cse | ({{13{FOR_I_and_4_cse}}, FOR_I_and_4_cse})
      | (signext_14_1(z_out_22[16])));
  assign memory_1_mux1h_10_nl = MUX1HOT_v_14_3_2((FOR_I_FOR_I_nor_1_nl), (BIAS_I_BIAS_I_nor_nl),
      (memory_2_rsci_q_d[14:1]), {memory_1_or_17_cse , memory_1_or_19_cse , (fsm_output[82])});
  assign memory_1_and_9_nl = MUX_v_14_2_2(14'b00000000000000, (memory_1_mux1h_10_nl),
      memory_1_or_seb);
  assign FOR_I_FOR_I_nor_2_nl = ~(FOR_I_nor_4_cse | FOR_I_and_4_cse);
  assign BIAS_I_BIAS_I_nor_3_nl = ~(FOR_I_nor_4_cse | (z_out_22[16]));
  assign memory_1_mux1h_11_nl = MUX1HOT_s_1_3_2((FOR_I_FOR_I_nor_2_nl), (BIAS_I_BIAS_I_nor_3_nl),
      (memory_2_rsci_q_d[0]), {memory_1_or_17_cse , memory_1_or_19_cse , (fsm_output[82])});
  assign memory_1_and_10_nl = (memory_1_mux1h_11_nl) & memory_1_or_seb;
  assign memory_1_rsci_d_d = {(memory_1_and_nl) , (memory_1_and_9_nl) , (memory_1_and_10_nl)};
  assign memory_1_rsci_we_d = or_dcpl_53 | (fsm_output[68]) | (fsm_output[55]) |
      (fsm_output[29]) | (fsm_output[3]) | (fsm_output[63]) | (fsm_output[42]) |
      (fsm_output[37]) | (fsm_output[16]) | (fsm_output[11]) | (fsm_output[82]);
  assign memory_1_rsci_re_d = (fsm_output[62]) | (fsm_output[36]) | (fsm_output[10])
      | (fsm_output[67]) | (fsm_output[41]) | (fsm_output[15]) | (fsm_output[87])
      | and_316_cse | and_317_cse | and_318_cse;
  assign nl_FOR_B_2_if_acc_12_nl = (FOR_B_2_if_acc_8_sdt_1[6:3]) + (CR2_simple_k_6_0_sva_5_0_1[3:0]);
  assign FOR_B_2_if_acc_12_nl = nl_FOR_B_2_if_acc_12_nl[3:0];
  assign nl_FOR_B_4_if_acc_16_nl = conv_s2u_4_6(FOR_B_4_if_acc_11_sdt_1[6:3]) + conv_u2u_5_6(CR3_simple_k_5_0_sva_4_0);
  assign FOR_B_4_if_acc_16_nl = nl_FOR_B_4_if_acc_16_nl[5:0];
  assign memory_2_mux1h_1_nl = MUX1HOT_v_8_3_2(({(FOR_B_2_if_acc_12_nl) , (FOR_B_2_if_acc_8_sdt_1[2:0])
      , (FOR_B_2_if_acc_9_psp_1[0])}), ({(FOR_B_4_if_acc_16_nl) , (FOR_B_4_if_acc_11_sdt_1[2:1])}),
      ({3'b0 , z_out_12}), {and_285_cse , and_283_cse , (fsm_output[81])});
  assign memory_2_not_4_nl = ~ memory_2_rsci_radr_d_mx0c0;
  assign memory_2_and_3_nl = MUX_v_8_2_2(8'b00000000, (memory_2_mux1h_1_nl), (memory_2_not_4_nl));
  assign memory_2_mux1h_4_nl = MUX1HOT_s_1_3_2((z_out_16[0]), (FOR_B_4_if_acc_11_sdt_1[0]),
      (z_out_11[2]), {and_285_cse , and_283_cse , (fsm_output[81])});
  assign memory_2_and_4_nl = (memory_2_mux1h_4_nl) & (~ memory_2_rsci_radr_d_mx0c0);
  assign memory_2_mux1h_5_nl = MUX1HOT_v_2_3_2((CR2_simple_j_aux_4_0_sva_1[1:0]),
      ({(FOR_B_4_if_acc_6_sdt_1[0]) , (CR3_simple_j_aux_3_0_sva_1[0])}), (z_out_11[1:0]),
      {and_285_cse , and_283_cse , (fsm_output[81])});
  assign memory_2_not_6_nl = ~ memory_2_rsci_radr_d_mx0c0;
  assign memory_2_and_5_nl = MUX_v_2_2_2(2'b00, (memory_2_mux1h_5_nl), (memory_2_not_6_nl));
  assign memory_2_rsci_radr_d = {(memory_2_and_3_nl) , (memory_2_and_4_nl) , (memory_2_and_5_nl)};
  assign nl_FOR_B_1_if_acc_5_nl = (FOR_B_1_if_acc_3_sdt_1[6:3]) + (MP1_simple_k_6_0_sva_5_0[3:0]);
  assign FOR_B_1_if_acc_5_nl = nl_FOR_B_1_if_acc_5_nl[3:0];
  assign nl_FOR_B_3_if_acc_5_nl = conv_u2u_3_6(z_out_10[5:3]) + conv_u2u_5_6(MP2_simple_k_5_0_sva_4_0);
  assign FOR_B_3_if_acc_5_nl = nl_FOR_B_3_if_acc_5_nl[5:0];
  assign memory_2_mux1h_nl = MUX1HOT_v_8_3_2(({(FOR_B_1_if_acc_5_nl) , (FOR_B_1_if_acc_3_sdt_1[2:0])
      , (z_out_23[0])}), ({(FOR_B_3_if_acc_5_nl) , (z_out_10[2:1])}), ({3'b0 , z_out_12}),
      {(fsm_output[24]) , (fsm_output[50]) , (fsm_output[76])});
  assign memory_2_not_1_nl = ~ memory_2_rsci_wadr_d_mx0c0;
  assign memory_2_and_nl = MUX_v_8_2_2(8'b00000000, (memory_2_mux1h_nl), (memory_2_not_1_nl));
  assign memory_2_mux1h_2_nl = MUX1HOT_s_1_3_2((z_out_8[0]), (z_out_10[0]), (z_out_21[2]),
      {(fsm_output[24]) , (fsm_output[50]) , (fsm_output[76])});
  assign memory_2_and_1_nl = (memory_2_mux1h_2_nl) & (~ memory_2_rsci_wadr_d_mx0c0);
  assign memory_2_mux1h_3_nl = MUX1HOT_v_2_3_2((MP1_simple_i_N_3_0_sva_1[1:0]), ({(FOR_B_3_if_acc_sdt_1[0])
      , (MP2_simple_i_N_2_0_sva_1[0])}), (z_out_21[1:0]), {(fsm_output[24]) , (fsm_output[50])
      , (fsm_output[76])});
  assign memory_2_not_3_nl = ~ memory_2_rsci_wadr_d_mx0c0;
  assign memory_2_and_2_nl = MUX_v_2_2_2(2'b00, (memory_2_mux1h_3_nl), (memory_2_not_3_nl));
  assign memory_2_rsci_wadr_d = {(memory_2_and_nl) , (memory_2_and_1_nl) , (memory_2_and_2_nl)};
  assign or_198_nl = (fsm_output[24]) | (fsm_output[0]);
  assign MP1_simple_bigger_mux1h_nl = MUX1HOT_v_16_3_2(MP1_simple_bigger_lpi_6_dfm_1,
      MP2_simple_bigger_lpi_6_dfm_1, MP3_simple_bigger_lpi_6_dfm_1, {(or_198_nl)
      , (fsm_output[50]) , (fsm_output[76])});
  assign memory_2_nand_nl = ~(and_dcpl_6 & (~ (fsm_output[24])) & (~ (fsm_output[0])));
  assign memory_2_rsci_d_d = MUX_v_16_2_2(16'b0000000000000000, (MP1_simple_bigger_mux1h_nl),
      (memory_2_nand_nl));
  assign memory_2_rsci_we_d = or_dcpl_53 | (fsm_output[76]) | (fsm_output[50]) |
      (fsm_output[24]);
  assign memory_2_rsci_re_d = and_283_cse | (fsm_output[81]) | and_285_cse;
  assign FOR_A_1_if_mux1h_4_cse = MUX1HOT_v_4_5_2(MP1_simple_j_4_1_sva, MP1_simple_j_N_3_0_sva_1,
      CR2_simple_i_1_3_0_sva, CR2_simple_i_2_3_0_sva, CR2_simple_i_3_0_sva, {(fsm_output[22])
      , (fsm_output[24]) , (fsm_output[29]) , (fsm_output[36]) , (fsm_output[41])});
  assign INIT_I_or_6_cse = (fsm_output[3]) | (fsm_output[10]) | (fsm_output[15]);
  assign INIT_I_or_4_cse = (fsm_output[74]) | (fsm_output[76]);
  always @(posedge clk) begin
    if ( rst ) begin
      reg_index_rsc_triosy_obj_ld_cse <= 1'b0;
      Prob_9_15_sva_2 <= 1'b0;
      Prob_9_0_sva_2 <= 1'b0;
      Prob_9_14_1_sva_2 <= 14'b0;
      Prob_8_15_sva_2 <= 1'b0;
      Prob_8_0_sva_2 <= 1'b0;
      Prob_8_14_1_sva_2 <= 14'b0;
      Prob_1_15_sva_2 <= 1'b0;
      Prob_1_0_sva_2 <= 1'b0;
      Prob_1_14_1_sva_2 <= 14'b0;
      Prob_7_15_sva_2 <= 1'b0;
      Prob_7_0_sva_2 <= 1'b0;
      Prob_7_14_1_sva_2 <= 14'b0;
      Prob_2_15_sva_2 <= 1'b0;
      Prob_2_0_sva_2 <= 1'b0;
      Prob_2_14_1_sva_2 <= 14'b0;
      Prob_6_15_sva_2 <= 1'b0;
      Prob_6_0_sva_2 <= 1'b0;
      Prob_6_14_1_sva_2 <= 14'b0;
      Prob_3_15_sva_2 <= 1'b0;
      Prob_3_0_sva_2 <= 1'b0;
      Prob_3_14_1_sva_2 <= 14'b0;
      Prob_5_15_sva_2 <= 1'b0;
      Prob_5_0_sva_2 <= 1'b0;
      Prob_5_14_1_sva_2 <= 14'b0;
      Prob_4_15_sva_2 <= 1'b0;
      Prob_4_0_sva_2 <= 1'b0;
      Prob_4_14_1_sva_2 <= 14'b0;
      CR1_simple_i_1_4_0_sva <= 5'b0;
      reg_INIT_I_slc_INIT_I_acc_2_cse <= 1'b0;
      CR1_simple_i_1_4_0_sva_1 <= 5'b0;
      CR1_simple_b_1_0_sva <= 2'b0;
      CR1_simple_b_1_0_sva_1 <= 2'b0;
      FOR_B_lor_2_lpi_7_dfm_st <= 1'b0;
      CR1_simple_aux_0_lpi_7_dfm <= 1'b0;
      CR1_simple_aux_14_1_lpi_7_dfm <= 14'b0;
      CR1_simple_aux_15_lpi_7_dfm <= 1'b0;
      reg_FOR_I_asn_CR1_simple_add_AF_10_FOR_I_acc_psp_cse <= 5'b0;
      CR1_simple_i_4_0_sva <= 5'b0;
      BIAS_I_slc_15_1_itm <= 15'b0;
      MP1_simple_j_N_3_0_sva <= 4'b0;
      MP1_simple_i_N_3_0_sva <= 4'b0;
      MP1_simple_a_1_0_sva <= 2'b0;
      reg_FOR_A_1_lor_lpi_6_dfm_cse <= 1'b0;
      CR2_simple_i_1_3_0_sva <= 4'b0;
      CR2_simple_i_1_3_0_sva_1 <= 4'b0;
      CR2_simple_b_1_0_sva <= 2'b0;
      FOR_B_2_lor_2_lpi_7_dfm_st <= 1'b0;
      CR2_simple_aux_0_lpi_7_dfm <= 1'b0;
      CR2_simple_aux_14_1_lpi_7_dfm <= 14'b0;
      CR2_simple_aux_15_lpi_7_dfm <= 1'b0;
      reg_FOR_I_2_acc_11_psp_cse <= 4'b0;
      reg_FOR_I_2_acc_9_sdt_cse <= 3'b0;
      reg_FOR_I_2_acc_10_psp_cse <= 1'b0;
      reg_FOR_I_2_acc_8_sdt_cse <= 1'b0;
      CR2_simple_i_3_0_sva <= 4'b0;
      BIAS_I_1_slc_15_1_itm <= 15'b0;
      MP2_simple_j_N_2_0_sva <= 3'b0;
      MP2_simple_i_N_2_0_sva <= 3'b0;
      MP2_simple_a_1_0_sva <= 2'b0;
      CR3_simple_i_1_2_0_sva <= 3'b0;
      CR3_simple_i_1_2_0_sva_1 <= 3'b0;
      CR3_simple_b_1_0_sva <= 2'b0;
      FOR_B_4_lor_2_lpi_7_dfm_st <= 1'b0;
      CR3_simple_aux_0_lpi_7_dfm <= 1'b0;
      CR3_simple_aux_14_1_lpi_7_dfm <= 14'b0;
      CR3_simple_aux_15_lpi_7_dfm <= 1'b0;
      reg_FOR_I_4_acc_11_psp_cse <= 5'b0;
      reg_FOR_I_4_acc_9_sdt_cse <= 3'b0;
      reg_FOR_I_4_acc_8_sdt_2_0_cse <= 1'b0;
      CR3_simple_i_2_0_sva <= 3'b0;
      BIAS_I_2_slc_15_1_itm <= 15'b0;
      MP3_simple_j_N_1_0_sva_1_1 <= 1'b0;
      MP3_simple_j_N_1_0_sva_0 <= 1'b0;
      MP3_simple_i_N_1_0_sva_1_1 <= 1'b0;
      MP3_simple_i_N_1_0_sva_0 <= 1'b0;
      reshape_simple_k_4_0_sva <= 5'b0;
      Prob_0_sva_2_15 <= 1'b0;
      Prob_0_sva_2_0 <= 1'b0;
      Prob_0_sva_2_14_1 <= 14'b0;
      perceptron_simple_k_7_0_sva <= 8'b0;
      FOR_K_7_slc_FOR_K_7_acc_6_itm <= 1'b0;
      FOR_K_7_mux_28_itm <= 1'b0;
      FOR_K_7_mux_29_itm <= 14'b0;
      FOR_K_7_mux_30_itm <= 1'b0;
      perceptron_simple_k_7_0_sva_1 <= 8'b0;
      k_sva <= 4'b0;
      max_sva_14_1 <= 14'b0;
      max_sva_15 <= 1'b0;
      max_sva_0 <= 1'b0;
    end
    else begin
      reg_index_rsc_triosy_obj_ld_cse <= (~ (z_out_7[3])) & (fsm_output[90]);
      Prob_9_15_sva_2 <= MUX_s_1_2_2((FOR_K_7_mux_1_nl), Prob_9_15_sva_2, or_tmp_125);
      Prob_9_0_sva_2 <= MUX_s_1_2_2((FOR_K_7_mux_2_nl), Prob_9_0_sva_2, or_tmp_125);
      Prob_9_14_1_sva_2 <= MUX1HOT_v_14_3_2(Prob_9_14_1_sva_1, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
          Prob_9_14_1_sva_2, {(Prob_Prob_nor_nl) , (Prob_and_19_nl) , or_tmp_125});
      Prob_8_15_sva_2 <= MUX_s_1_2_2((FOR_K_7_mux_4_nl), Prob_8_15_sva_2, or_tmp_125);
      Prob_8_0_sva_2 <= MUX_s_1_2_2((FOR_K_7_mux_5_nl), Prob_8_0_sva_2, or_tmp_125);
      Prob_8_14_1_sva_2 <= MUX1HOT_v_14_3_2(Prob_8_14_1_sva_1, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
          Prob_8_14_1_sva_2, {(Prob_Prob_nor_1_nl) , (Prob_and_17_nl) , or_tmp_125});
      Prob_1_15_sva_2 <= MUX_s_1_2_2((FOR_K_7_mux_7_nl), Prob_1_15_sva_2, or_tmp_125);
      Prob_1_0_sva_2 <= MUX_s_1_2_2((FOR_K_7_mux_8_nl), Prob_1_0_sva_2, or_tmp_125);
      Prob_1_14_1_sva_2 <= MUX1HOT_v_14_3_2(Prob_1_14_1_sva_1, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
          Prob_1_14_1_sva_2, {(Prob_Prob_nor_2_nl) , (Prob_and_15_nl) , or_tmp_125});
      Prob_7_15_sva_2 <= MUX_s_1_2_2((FOR_K_7_mux_10_nl), Prob_7_15_sva_2, or_tmp_125);
      Prob_7_0_sva_2 <= MUX_s_1_2_2((FOR_K_7_mux_11_nl), Prob_7_0_sva_2, or_tmp_125);
      Prob_7_14_1_sva_2 <= MUX1HOT_v_14_3_2(Prob_7_14_1_sva_1, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
          Prob_7_14_1_sva_2, {(Prob_Prob_nor_3_nl) , (Prob_and_13_nl) , or_tmp_125});
      Prob_2_15_sva_2 <= MUX_s_1_2_2((FOR_K_7_mux_13_nl), Prob_2_15_sva_2, or_tmp_125);
      Prob_2_0_sva_2 <= MUX_s_1_2_2((FOR_K_7_mux_14_nl), Prob_2_0_sva_2, or_tmp_125);
      Prob_2_14_1_sva_2 <= MUX1HOT_v_14_3_2(Prob_2_14_1_sva_1, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
          Prob_2_14_1_sva_2, {(Prob_Prob_nor_4_nl) , (Prob_and_11_nl) , or_tmp_125});
      Prob_6_15_sva_2 <= MUX_s_1_2_2((FOR_K_7_mux_16_nl), Prob_6_15_sva_2, or_tmp_125);
      Prob_6_0_sva_2 <= MUX_s_1_2_2((FOR_K_7_mux_17_nl), Prob_6_0_sva_2, or_tmp_125);
      Prob_6_14_1_sva_2 <= MUX1HOT_v_14_3_2(Prob_6_14_1_sva_1, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
          Prob_6_14_1_sva_2, {(Prob_Prob_nor_5_nl) , (Prob_and_9_nl) , or_tmp_125});
      Prob_3_15_sva_2 <= MUX_s_1_2_2((FOR_K_7_mux_19_nl), Prob_3_15_sva_2, or_tmp_125);
      Prob_3_0_sva_2 <= MUX_s_1_2_2((FOR_K_7_mux_20_nl), Prob_3_0_sva_2, or_tmp_125);
      Prob_3_14_1_sva_2 <= MUX1HOT_v_14_3_2(Prob_3_14_1_sva_1, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
          Prob_3_14_1_sva_2, {(Prob_Prob_nor_6_nl) , (Prob_and_7_nl) , or_tmp_125});
      Prob_5_15_sva_2 <= MUX_s_1_2_2((FOR_K_7_mux_22_nl), Prob_5_15_sva_2, or_tmp_125);
      Prob_5_0_sva_2 <= MUX_s_1_2_2((FOR_K_7_mux_23_nl), Prob_5_0_sva_2, or_tmp_125);
      Prob_5_14_1_sva_2 <= MUX1HOT_v_14_3_2(Prob_5_14_1_sva_1, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
          Prob_5_14_1_sva_2, {(Prob_Prob_nor_7_nl) , (Prob_and_5_nl) , or_tmp_125});
      Prob_4_15_sva_2 <= MUX_s_1_2_2((FOR_K_7_mux_25_nl), Prob_4_15_sva_2, or_tmp_125);
      Prob_4_0_sva_2 <= MUX_s_1_2_2((FOR_K_7_mux_26_nl), Prob_4_0_sva_2, or_tmp_125);
      Prob_4_14_1_sva_2 <= MUX1HOT_v_14_3_2(Prob_4_14_1_sva_1, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
          Prob_4_14_1_sva_2, {(Prob_Prob_nor_8_nl) , (Prob_and_3_nl) , or_tmp_125});
      CR1_simple_i_1_4_0_sva <= MUX_v_5_2_2(5'b00000, CR1_simple_i_1_4_0_sva_1, (CR1_simple_i_nor_nl));
      reg_INIT_I_slc_INIT_I_acc_2_cse <= z_out[2];
      CR1_simple_i_1_4_0_sva_1 <= z_out_9;
      CR1_simple_b_1_0_sva <= MUX_v_2_2_2(2'b00, CR1_simple_b_1_0_sva_1, (fsm_output[8]));
      CR1_simple_b_1_0_sva_1 <= z_out_2[1:0];
      FOR_B_lor_2_lpi_7_dfm_st <= or_125_cse;
      CR1_simple_aux_0_lpi_7_dfm <= MUX_s_1_2_2(CR1_simple_aux_0_lpi_7_mx1, CR1_simple_aux_0_lpi_7_dfm,
          and_4_cse);
      CR1_simple_aux_14_1_lpi_7_dfm <= MUX_v_14_2_2(CR1_simple_aux_14_1_lpi_7_mx1,
          CR1_simple_aux_14_1_lpi_7_dfm, and_4_cse);
      CR1_simple_aux_15_lpi_7_dfm <= MUX_s_1_2_2(CR1_simple_aux_15_lpi_7_mx1, CR1_simple_aux_15_lpi_7_dfm,
          and_4_cse);
      reg_FOR_I_asn_CR1_simple_add_AF_10_FOR_I_acc_psp_cse <= z_out_19;
      CR1_simple_i_4_0_sva <= MUX_v_5_2_2(5'b00000, CR1_simple_i_4_0_sva_1, (fsm_output[17]));
      BIAS_I_slc_15_1_itm <= B_1_rsci_q_d[15:1];
      MP1_simple_j_N_3_0_sva <= MUX_v_4_2_2(MP1_simple_j_N_3_0_sva_1, 4'b1111, (not_408_nl));
      MP1_simple_i_N_3_0_sva <= MUX_v_4_2_2(MP1_simple_i_N_3_0_sva_1, 4'b1111, (MP1_simple_i_N_not_nl));
      MP1_simple_a_1_0_sva <= MUX_v_2_2_2(2'b00, CR1_simple_b_1_0_sva_1, (MP1_simple_a_nor_nl));
      reg_FOR_A_1_lor_lpi_6_dfm_cse <= nand_cse_1;
      CR2_simple_i_1_3_0_sva <= MUX_v_4_2_2(4'b0000, CR2_simple_i_1_3_0_sva_1, (fsm_output[30]));
      CR2_simple_i_1_3_0_sva_1 <= z_out_5;
      CR2_simple_b_1_0_sva <= MUX_v_2_2_2(2'b00, CR1_simple_b_1_0_sva_1, (fsm_output[34]));
      FOR_B_2_lor_2_lpi_7_dfm_st <= FOR_B_2_if_FOR_B_2_if_or_cse;
      CR2_simple_aux_0_lpi_7_dfm <= MUX_s_1_2_2(CR2_simple_aux_0_lpi_7_mx1, CR2_simple_aux_0_lpi_7_dfm,
          and_10_cse);
      CR2_simple_aux_14_1_lpi_7_dfm <= MUX_v_14_2_2(CR2_simple_aux_14_1_lpi_7_mx1,
          CR2_simple_aux_14_1_lpi_7_dfm, and_10_cse);
      CR2_simple_aux_15_lpi_7_dfm <= MUX_s_1_2_2(CR2_simple_aux_15_lpi_7_mx1, CR2_simple_aux_15_lpi_7_dfm,
          and_10_cse);
      reg_FOR_I_2_acc_11_psp_cse <= z_out_7;
      reg_FOR_I_2_acc_9_sdt_cse <= z_out_10[2:0];
      reg_FOR_I_2_acc_10_psp_cse <= z_out_23[0];
      reg_FOR_I_2_acc_8_sdt_cse <= z_out_8[0];
      CR2_simple_i_3_0_sva <= MUX_v_4_2_2(4'b0000, CR2_simple_i_3_0_sva_1, (fsm_output[43]));
      BIAS_I_1_slc_15_1_itm <= B_2_rsci_q_d[15:1];
      MP2_simple_j_N_2_0_sva <= MUX_v_3_2_2(MP2_simple_j_N_2_0_sva_1, 3'b111, (not_404_nl));
      MP2_simple_i_N_2_0_sva <= MUX_v_3_2_2(MP2_simple_i_N_2_0_sva_1, 3'b111, (MP2_simple_i_N_not_nl));
      MP2_simple_a_1_0_sva <= MUX_v_2_2_2(2'b00, CR1_simple_b_1_0_sva_1, (MP2_simple_a_nor_nl));
      CR3_simple_i_1_2_0_sva <= MUX_v_3_2_2(3'b000, CR3_simple_i_1_2_0_sva_1, (fsm_output[56]));
      CR3_simple_i_1_2_0_sva_1 <= z_out_6;
      CR3_simple_b_1_0_sva <= MUX_v_2_2_2(2'b00, CR1_simple_b_1_0_sva_1, (fsm_output[60]));
      FOR_B_4_lor_2_lpi_7_dfm_st <= FOR_B_4_if_FOR_B_4_if_or_cse;
      CR3_simple_aux_0_lpi_7_dfm <= MUX_s_1_2_2(CR3_simple_aux_0_lpi_7_mx1, CR3_simple_aux_0_lpi_7_dfm,
          and_16_cse);
      CR3_simple_aux_14_1_lpi_7_dfm <= MUX_v_14_2_2(CR3_simple_aux_14_1_lpi_7_mx1,
          CR3_simple_aux_14_1_lpi_7_dfm, and_16_cse);
      CR3_simple_aux_15_lpi_7_dfm <= MUX_s_1_2_2(CR3_simple_aux_15_lpi_7_mx1, CR3_simple_aux_15_lpi_7_dfm,
          and_16_cse);
      reg_FOR_I_4_acc_11_psp_cse <= z_out_12;
      reg_FOR_I_4_acc_9_sdt_cse <= z_out_20[2:0];
      reg_FOR_I_4_acc_8_sdt_2_0_cse <= z_out_27_2_0[0];
      CR3_simple_i_2_0_sva <= MUX_v_3_2_2(3'b000, CR3_simple_i_2_0_sva_1, (fsm_output[69]));
      BIAS_I_2_slc_15_1_itm <= B_3_rsci_q_d[15:1];
      MP3_simple_j_N_1_0_sva_1_1 <= ~ (fsm_output[79]);
      MP3_simple_j_N_1_0_sva_0 <= (MP3_simple_j_N_1_0_sva_1[0]) | (~ (fsm_output[79]));
      MP3_simple_i_N_1_0_sva_1_1 <= ~ (fsm_output[78]);
      MP3_simple_i_N_1_0_sva_0 <= (MP3_simple_i_N_1_0_sva_1[0]) | (~ (fsm_output[78]));
      reshape_simple_k_4_0_sva <= MUX_v_5_2_2(5'b00000, reshape_simple_k_4_0_sva_1,
          (fsm_output[83]));
      Prob_0_sva_2_15 <= MUX_s_1_2_2((FOR_K_7_mux_28_nl), Prob_0_sva_2_15, or_tmp_376);
      Prob_0_sva_2_0 <= MUX_s_1_2_2((FOR_K_7_mux_29_nl), Prob_0_sva_2_0, or_tmp_376);
      Prob_0_sva_2_14_1 <= MUX1HOT_v_14_3_2(Prob_0_sva_1_14_1, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
          Prob_0_sva_2_14_1, {(Prob_Prob_nor_9_nl) , (Prob_and_1_nl) , or_tmp_376});
      perceptron_simple_k_7_0_sva <= MUX_v_8_2_2(8'b00000000, perceptron_simple_k_7_0_sva_1,
          (fsm_output[88]));
      FOR_K_7_slc_FOR_K_7_acc_6_itm <= readslicef_7_1_6((FOR_K_7_acc_nl));
      FOR_K_7_mux_28_itm <= MUX_s_1_10_2(Prob_0_sva_1_15, Prob_1_15_sva_1, Prob_2_15_sva_1,
          Prob_3_15_sva_1, Prob_4_15_sva_1, Prob_5_15_sva_1, Prob_6_15_sva_1, Prob_7_15_sva_1,
          Prob_8_15_sva_1, Prob_9_15_sva_1, perceptron_simple_j_3_0_sva);
      FOR_K_7_mux_29_itm <= MUX_v_14_10_2(Prob_0_sva_1_14_1, Prob_1_14_1_sva_1, Prob_2_14_1_sva_1,
          Prob_3_14_1_sva_1, Prob_4_14_1_sva_1, Prob_5_14_1_sva_1, Prob_6_14_1_sva_1,
          Prob_7_14_1_sva_1, Prob_8_14_1_sva_1, Prob_9_14_1_sva_1, perceptron_simple_j_3_0_sva);
      FOR_K_7_mux_30_itm <= MUX_s_1_10_2(Prob_0_sva_1_0, Prob_1_0_sva_1, Prob_2_0_sva_1,
          Prob_3_0_sva_1, Prob_4_0_sva_1, Prob_5_0_sva_1, Prob_6_0_sva_1, Prob_7_0_sva_1,
          Prob_8_0_sva_1, Prob_9_0_sva_1, perceptron_simple_j_3_0_sva);
      perceptron_simple_k_7_0_sva_1 <= perceptron_simple_k_7_0_sva_2;
      k_sva <= MUX_v_4_2_2(4'b0000, z_out_5, (fsm_output[90]));
      max_sva_14_1 <= MUX_v_14_2_2(Prob_0_sva_2_14_1, max_sva_14_1_mx1, fsm_output[90]);
      max_sva_15 <= MUX_s_1_2_2(Prob_0_sva_2_15, (for_mux_1_nl), fsm_output[90]);
      max_sva_0 <= MUX_s_1_2_2(Prob_0_sva_2_0, (for_mux_2_nl), fsm_output[90]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      index_rsci_idat <= 4'b0;
    end
    else if ( ~((~ (fsm_output[90])) | (z_out_7[3])) ) begin
      index_rsci_idat <= max_sva_14_1_mx1[10:7];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR1_simple_l_1_6_0_sva_5_0 <= 6'b0;
    end
    else if ( reg_CR1_simple_l_1_6_0_sva_5_CR1_simple_l_or_cse ) begin
      CR1_simple_l_1_6_0_sva_5_0 <= MUX_v_6_2_2(6'b000000, (z_out_13[5:0]), (CR1_simple_l_not_1_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR1_simple_j_1_4_0_sva <= 5'b0;
    end
    else if ( (fsm_output[5]) | reg_CR1_simple_l_1_6_0_sva_5_CR1_simple_l_or_cse
        ) begin
      CR1_simple_j_1_4_0_sva <= MUX_v_5_2_2(5'b00000, z_out_9, (CR1_simple_j_not_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR1_simple_k_1_0_sva <= 2'b0;
    end
    else if ( (fsm_output[19]) | (fsm_output[6]) | (fsm_output[14]) ) begin
      CR1_simple_k_1_0_sva <= MUX_v_2_2_2(2'b00, (z_out_2[1:0]), (fsm_output[14]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR1_simple_a_1_0_sva <= 2'b0;
    end
    else if ( or_332_cse | (fsm_output[9]) ) begin
      CR1_simple_a_1_0_sva <= MUX_v_2_2_2(2'b00, (z_out_2[1:0]), (fsm_output[9]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR1_simple_l_6_0_sva_5_0_1 <= 6'b0;
    end
    else if ( (fsm_output[6]) | (fsm_output[19]) ) begin
      CR1_simple_l_6_0_sva_5_0_1 <= MUX_v_6_2_2(6'b000000, (z_out_13[5:0]), (fsm_output[19]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR1_simple_aux_15_lpi_7 <= 1'b0;
      CR1_simple_aux_14_1_lpi_7 <= 14'b0;
      CR1_simple_aux_0_lpi_7 <= 1'b0;
    end
    else if ( reg_CR1_simple_CR1_simple_aux_or_1_cse ) begin
      CR1_simple_aux_15_lpi_7 <= (CR1_simple_aux_mux_14_nl) & (~ or_332_cse);
      CR1_simple_aux_14_1_lpi_7 <= MUX_v_14_2_2(14'b00000000000000, (CR1_simple_aux_mux_13_nl),
          (not_410_nl));
      CR1_simple_aux_0_lpi_7 <= (CR1_simple_aux_mux_12_nl) & (~ or_332_cse);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR1_simple_j_2_4_0_sva <= 5'b0;
    end
    else if ( (fsm_output[19]) | (fsm_output[14]) | (fsm_output[6]) | (fsm_output[13])
        ) begin
      CR1_simple_j_2_4_0_sva <= MUX_v_5_2_2(5'b00000, z_out_9, (fsm_output[13]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR1_simple_i_2_4_0_sva <= 5'b0;
    end
    else if ( or_332_cse ) begin
      CR1_simple_i_2_4_0_sva <= MUX_v_5_2_2(5'b00000, CR1_simple_i_2_4_0_sva_1, (fsm_output[12]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      FOR_I_slc_FOR_I_acc_2_itm <= 1'b0;
    end
    else if ( fsm_output[10] ) begin
      FOR_I_slc_FOR_I_acc_2_itm <= z_out[2];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR1_simple_i_2_4_0_sva_1 <= 5'b0;
    end
    else if ( fsm_output[10] ) begin
      CR1_simple_i_2_4_0_sva_1 <= z_out_9;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR1_simple_j_4_0_sva <= 5'b0;
    end
    else if ( (fsm_output[14]) | (fsm_output[18]) ) begin
      CR1_simple_j_4_0_sva <= MUX_v_5_2_2(5'b00000, z_out_9, (fsm_output[18]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      BIAS_I_slc_BIAS_I_acc_2_itm <= 1'b0;
    end
    else if ( fsm_output[15] ) begin
      BIAS_I_slc_BIAS_I_acc_2_itm <= z_out[2];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR1_simple_i_4_0_sva_1 <= 5'b0;
    end
    else if ( fsm_output[15] ) begin
      CR1_simple_i_4_0_sva_1 <= z_out_9;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP1_simple_k_6_0_sva_5_0 <= 6'b0;
    end
    else if ( (fsm_output[19]) | (fsm_output[28]) ) begin
      MP1_simple_k_6_0_sva_5_0 <= MUX_v_6_2_2(6'b000000, (z_out_13[5:0]), (fsm_output[28]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP1_simple_j_4_1_sva <= 4'b0;
    end
    else if ( (fsm_output[28]) | (fsm_output[19]) | (fsm_output[27]) ) begin
      MP1_simple_j_4_1_sva <= MUX_v_4_2_2(4'b0000, z_out_5, (fsm_output[27]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP1_simple_i_4_1_sva <= 4'b0;
    end
    else if ( (fsm_output[20]) | (fsm_output[26]) ) begin
      MP1_simple_i_4_1_sva <= MUX_v_4_2_2(4'b0000, z_out_5, (MP1_simple_i_not_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP1_simple_j_N_3_0_sva_1 <= 4'b0;
    end
    else if ( fsm_output[20] ) begin
      MP1_simple_j_N_3_0_sva_1 <= z_out_5;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP1_simple_b_1_0_sva <= 2'b0;
    end
    else if ( (fsm_output[21]) | (fsm_output[25]) ) begin
      MP1_simple_b_1_0_sva <= MUX_v_2_2_2(2'b00, CR1_simple_b_1_0_sva_1, (MP1_simple_b_not_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP1_simple_bigger_lpi_6 <= 16'b0;
    end
    else if ( (fsm_output[21]) | (fsm_output[23]) | (fsm_output[25]) ) begin
      MP1_simple_bigger_lpi_6 <= MUX_v_16_2_2(16'b0000000000000000, (memory_1_mux_3_nl),
          (MP1_simple_bigger_not_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP1_simple_i_N_3_0_sva_1 <= 4'b0;
    end
    else if ( fsm_output[21] ) begin
      MP1_simple_i_N_3_0_sva_1 <= z_out_5;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP1_simple_bigger_lpi_6_dfm_1 <= 16'b0;
    end
    else if ( fsm_output[23] ) begin
      MP1_simple_bigger_lpi_6_dfm_1 <= MP1_simple_bigger_lpi_6_mx1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR2_simple_l_1_5_0_sva_4_0 <= 5'b0;
    end
    else if ( (fsm_output[28]) | (fsm_output[32]) ) begin
      CR2_simple_l_1_5_0_sva_4_0 <= MUX_v_5_2_2(5'b00000, (z_out_16[4:0]), (fsm_output[32]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR2_simple_j_1_3_0_sva <= 4'b0;
    end
    else if ( (fsm_output[32]) | (fsm_output[28]) | (fsm_output[31]) ) begin
      CR2_simple_j_1_3_0_sva <= MUX_v_4_2_2(4'b0000, z_out_5, (fsm_output[31]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR2_simple_k_6_0_sva_5_0_1 <= 6'b0;
    end
    else if ( (fsm_output[45]) | (fsm_output[32]) | (fsm_output[40]) ) begin
      CR2_simple_k_6_0_sva_5_0_1 <= MUX_v_6_2_2(6'b000000, (z_out_13[5:0]), (fsm_output[40]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR2_simple_a_1_0_sva <= 2'b0;
    end
    else if ( or_400_cse | (fsm_output[35]) ) begin
      CR2_simple_a_1_0_sva <= MUX_v_2_2_2(2'b00, (z_out_2[1:0]), (fsm_output[35]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR2_simple_l_5_0_sva_4_0_1 <= 5'b0;
    end
    else if ( (fsm_output[32]) | (fsm_output[45]) ) begin
      CR2_simple_l_5_0_sva_4_0_1 <= MUX_v_5_2_2(5'b00000, (z_out_16[4:0]), (fsm_output[45]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR2_simple_aux_15_lpi_7 <= 1'b0;
      CR2_simple_aux_14_1_lpi_7 <= 14'b0;
      CR2_simple_aux_0_lpi_7 <= 1'b0;
    end
    else if ( reg_CR2_simple_CR2_simple_aux_or_1_cse ) begin
      CR2_simple_aux_15_lpi_7 <= (CR1_simple_aux_mux_11_nl) & (~ or_400_cse);
      CR2_simple_aux_14_1_lpi_7 <= MUX_v_14_2_2(14'b00000000000000, (CR1_simple_aux_mux_10_nl),
          (not_406_nl));
      CR2_simple_aux_0_lpi_7 <= (CR1_simple_aux_mux_9_nl) & (~ or_400_cse);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR2_simple_j_2_3_0_sva <= 4'b0;
    end
    else if ( (fsm_output[45]) | (fsm_output[40]) | (fsm_output[32]) | (fsm_output[39])
        ) begin
      CR2_simple_j_2_3_0_sva <= MUX_v_4_2_2(4'b0000, z_out_5, (fsm_output[39]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR2_simple_i_2_3_0_sva <= 4'b0;
    end
    else if ( or_400_cse ) begin
      CR2_simple_i_2_3_0_sva <= MUX_v_4_2_2(4'b0000, CR2_simple_i_2_3_0_sva_1, (fsm_output[38]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      FOR_I_2_slc_FOR_I_2_acc_2_itm <= 1'b0;
    end
    else if ( fsm_output[36] ) begin
      FOR_I_2_slc_FOR_I_2_acc_2_itm <= z_out[2];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR2_simple_i_2_3_0_sva_1 <= 4'b0;
    end
    else if ( fsm_output[36] ) begin
      CR2_simple_i_2_3_0_sva_1 <= z_out_5;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR2_simple_j_3_0_sva <= 4'b0;
    end
    else if ( (fsm_output[40]) | (fsm_output[44]) ) begin
      CR2_simple_j_3_0_sva <= MUX_v_4_2_2(4'b0000, z_out_5, (fsm_output[44]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      BIAS_I_1_slc_BIAS_I_1_acc_2_itm <= 1'b0;
    end
    else if ( fsm_output[41] ) begin
      BIAS_I_1_slc_BIAS_I_1_acc_2_itm <= z_out[2];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR2_simple_i_3_0_sva_1 <= 4'b0;
    end
    else if ( fsm_output[41] ) begin
      CR2_simple_i_3_0_sva_1 <= z_out_5;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP2_simple_k_5_0_sva_4_0 <= 5'b0;
    end
    else if ( (fsm_output[45]) | (fsm_output[54]) ) begin
      MP2_simple_k_5_0_sva_4_0 <= MUX_v_5_2_2(5'b00000, (z_out_16[4:0]), (fsm_output[54]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP2_simple_j_3_1_sva <= 3'b0;
    end
    else if ( (fsm_output[54]) | (fsm_output[45]) | (fsm_output[53]) ) begin
      MP2_simple_j_3_1_sva <= MUX_v_3_2_2(3'b000, z_out_6, (fsm_output[53]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP2_simple_i_3_1_sva <= 3'b0;
    end
    else if ( (fsm_output[46]) | (fsm_output[52]) ) begin
      MP2_simple_i_3_1_sva <= MUX_v_3_2_2(3'b000, z_out_6, (MP2_simple_i_not_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP2_simple_j_N_2_0_sva_1 <= 3'b0;
    end
    else if ( fsm_output[46] ) begin
      MP2_simple_j_N_2_0_sva_1 <= z_out_6;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP2_simple_b_1_0_sva <= 2'b0;
    end
    else if ( (fsm_output[47]) | (fsm_output[51]) ) begin
      MP2_simple_b_1_0_sva <= MUX_v_2_2_2(2'b00, CR1_simple_b_1_0_sva_1, (MP2_simple_b_not_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP2_simple_bigger_lpi_6 <= 16'b0;
    end
    else if ( (fsm_output[47]) | (fsm_output[49]) | (fsm_output[51]) ) begin
      MP2_simple_bigger_lpi_6 <= MUX_v_16_2_2(16'b0000000000000000, (memory_1_mux_4_nl),
          (MP2_simple_bigger_not_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP2_simple_i_N_2_0_sva_1 <= 3'b0;
    end
    else if ( fsm_output[47] ) begin
      MP2_simple_i_N_2_0_sva_1 <= z_out_6;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP2_simple_bigger_lpi_6_dfm_1 <= 16'b0;
    end
    else if ( fsm_output[49] ) begin
      MP2_simple_bigger_lpi_6_dfm_1 <= MP2_simple_bigger_lpi_6_mx1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR3_simple_l_1_4_0_sva <= 5'b0;
    end
    else if ( (fsm_output[54]) | (fsm_output[58]) ) begin
      CR3_simple_l_1_4_0_sva <= MUX_v_5_2_2(5'b00000, z_out_9, (fsm_output[58]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR3_simple_j_1_2_0_sva <= 3'b0;
    end
    else if ( (fsm_output[58]) | (fsm_output[54]) | (fsm_output[57]) ) begin
      CR3_simple_j_1_2_0_sva <= MUX_v_3_2_2(3'b000, z_out_6, (fsm_output[57]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR3_simple_k_5_0_sva_4_0 <= 5'b0;
    end
    else if ( (fsm_output[71]) | (fsm_output[58]) | (fsm_output[66]) ) begin
      CR3_simple_k_5_0_sva_4_0 <= MUX_v_5_2_2(5'b00000, (z_out_16[4:0]), (fsm_output[66]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR3_simple_a_1_0_sva <= 2'b0;
    end
    else if ( or_468_cse | (fsm_output[61]) ) begin
      CR3_simple_a_1_0_sva <= MUX_v_2_2_2(2'b00, (z_out_2[1:0]), (fsm_output[61]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR3_simple_l_4_0_sva <= 5'b0;
    end
    else if ( (fsm_output[58]) | (fsm_output[71]) ) begin
      CR3_simple_l_4_0_sva <= MUX_v_5_2_2(5'b00000, z_out_9, (fsm_output[71]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR3_simple_aux_15_lpi_7 <= 1'b0;
      CR3_simple_aux_14_1_lpi_7 <= 14'b0;
      CR3_simple_aux_0_lpi_7 <= 1'b0;
    end
    else if ( reg_CR3_simple_CR3_simple_aux_or_1_cse ) begin
      CR3_simple_aux_15_lpi_7 <= (CR1_simple_aux_mux_8_nl) & (~ or_468_cse);
      CR3_simple_aux_14_1_lpi_7 <= MUX_v_14_2_2(14'b00000000000000, (CR1_simple_aux_mux_7_nl),
          (not_402_nl));
      CR3_simple_aux_0_lpi_7 <= (CR1_simple_aux_mux_6_nl) & (~ or_468_cse);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR3_simple_j_2_2_0_sva <= 3'b0;
    end
    else if ( (fsm_output[71]) | (fsm_output[66]) | (fsm_output[58]) | (fsm_output[65])
        ) begin
      CR3_simple_j_2_2_0_sva <= MUX_v_3_2_2(3'b000, z_out_6, (fsm_output[65]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR3_simple_i_2_2_0_sva <= 3'b0;
    end
    else if ( or_468_cse ) begin
      CR3_simple_i_2_2_0_sva <= MUX_v_3_2_2(3'b000, CR3_simple_i_2_2_0_sva_1, (fsm_output[64]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      FOR_I_4_slc_FOR_I_4_acc_2_itm <= 1'b0;
    end
    else if ( fsm_output[62] ) begin
      FOR_I_4_slc_FOR_I_4_acc_2_itm <= z_out[2];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR3_simple_i_2_2_0_sva_1 <= 3'b0;
    end
    else if ( fsm_output[62] ) begin
      CR3_simple_i_2_2_0_sva_1 <= z_out_6;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR3_simple_j_2_0_sva <= 3'b0;
    end
    else if ( (fsm_output[66]) | (fsm_output[70]) ) begin
      CR3_simple_j_2_0_sva <= MUX_v_3_2_2(3'b000, z_out_6, (fsm_output[70]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      BIAS_I_2_slc_BIAS_I_2_acc_2_itm <= 1'b0;
    end
    else if ( fsm_output[67] ) begin
      BIAS_I_2_slc_BIAS_I_2_acc_2_itm <= z_out[2];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      CR3_simple_i_2_0_sva_1 <= 3'b0;
    end
    else if ( fsm_output[67] ) begin
      CR3_simple_i_2_0_sva_1 <= z_out_6;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP3_simple_k_4_0_sva <= 5'b0;
    end
    else if ( (fsm_output[71]) | (fsm_output[80]) ) begin
      MP3_simple_k_4_0_sva <= MUX_v_5_2_2(5'b00000, z_out_9, (fsm_output[80]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP3_simple_j_2_1_sva <= 2'b0;
    end
    else if ( (fsm_output[71]) | (fsm_output[80]) | (fsm_output[79]) ) begin
      MP3_simple_j_2_1_sva <= MUX_v_2_2_2(2'b00, (z_out_2[1:0]), (fsm_output[79]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP3_simple_i_2_1_sva <= 2'b0;
    end
    else if ( (fsm_output[72]) | (fsm_output[78]) ) begin
      MP3_simple_i_2_1_sva <= MUX_v_2_2_2(2'b00, (z_out_2[1:0]), (MP3_simple_i_not_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP3_simple_j_N_1_0_sva_1 <= 2'b0;
    end
    else if ( fsm_output[72] ) begin
      MP3_simple_j_N_1_0_sva_1 <= z_out_2[1:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP3_simple_a_1_0_sva <= 2'b0;
    end
    else if ( (fsm_output[75]) | reg_MP3_simple_b_1_MP3_simple_b_or_cse ) begin
      MP3_simple_a_1_0_sva <= MUX_v_2_2_2(2'b00, CR1_simple_b_1_0_sva_1, (MP3_simple_a_not_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP3_simple_b_1_0_sva <= 2'b0;
    end
    else if ( reg_MP3_simple_b_1_MP3_simple_b_or_cse ) begin
      MP3_simple_b_1_0_sva <= MUX_v_2_2_2(2'b00, CR1_simple_b_1_0_sva_1, (MP3_simple_b_not_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP3_simple_bigger_lpi_6 <= 16'b0;
    end
    else if ( (fsm_output[73]) | (fsm_output[75]) | (fsm_output[77]) ) begin
      MP3_simple_bigger_lpi_6 <= MUX_v_16_2_2(16'b0000000000000000, (memory_1_mux_5_nl),
          (MP3_simple_bigger_not_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP3_simple_i_N_1_0_sva_1 <= 2'b0;
    end
    else if ( fsm_output[73] ) begin
      MP3_simple_i_N_1_0_sva_1 <= z_out_2[1:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MP3_simple_bigger_lpi_6_dfm_1 <= 16'b0;
    end
    else if ( fsm_output[75] ) begin
      MP3_simple_bigger_lpi_6_dfm_1 <= MP3_simple_bigger_lpi_6_mx1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reshape_simple_i_1_0_sva <= 2'b0;
    end
    else if ( (fsm_output[80]) | (fsm_output[85]) ) begin
      reshape_simple_i_1_0_sva <= MUX_v_2_2_2(2'b00, (z_out_2[1:0]), (fsm_output[85]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reshape_simple_j_1_0_sva <= 2'b0;
    end
    else if ( (fsm_output[85]) | (fsm_output[80]) | (fsm_output[84]) ) begin
      reshape_simple_j_1_0_sva <= MUX_v_2_2_2(2'b00, (z_out_2[1:0]), (fsm_output[84]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reshape_simple_add_N_10_0_lpi_4 <= 11'b0;
    end
    else if ( (fsm_output[80]) | reshape_simple_add_N_10_0_lpi_4_mx0c1 ) begin
      reshape_simple_add_N_10_0_lpi_4 <= MUX_v_11_2_2(11'b00000000000, reshape_simple_add_N_10_0_sva_1,
          reshape_simple_add_N_10_0_lpi_4_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      FOR_K_6_slc_FOR_K_6_acc_3_itm <= 1'b0;
    end
    else if ( fsm_output[81] ) begin
      FOR_K_6_slc_FOR_K_6_acc_3_itm <= z_out_7[3];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reshape_simple_k_4_0_sva_1 <= 5'b0;
    end
    else if ( fsm_output[81] ) begin
      reshape_simple_k_4_0_sva_1 <= z_out_9;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reshape_simple_add_N_10_0_sva_1 <= 11'b0;
    end
    else if ( ~((fsm_output[84:82]!=3'b000)) ) begin
      reshape_simple_add_N_10_0_sva_1 <= nl_reshape_simple_add_N_10_0_sva_1[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      perceptron_simple_j_3_0_sva <= 4'b0;
    end
    else if ( (fsm_output[85]) | (fsm_output[89]) ) begin
      perceptron_simple_j_3_0_sva <= MUX_v_4_2_2(4'b0000, z_out_5, (fsm_output[89]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_9_15_sva_1 <= 1'b0;
    end
    else if ( ~ FOR_J_7_or_29_rgt ) begin
      Prob_9_15_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d[15]), Prob_9_15_sva_2, (FOR_K_7_acc_7_psp_sva_1[16]),
          {or_tmp_379 , or_tmp_380 , FOR_J_7_and_81_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      FOR_J_7_and_21_cse_sva <= 1'b0;
    end
    else if ( ~ or_tmp_383 ) begin
      FOR_J_7_and_21_cse_sva <= FOR_J_7_and_stg_2_1_sva_1 & (perceptron_simple_j_3_0_sva[3]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_9_0_sva_1 <= 1'b0;
    end
    else if ( ~ FOR_J_7_or_29_rgt ) begin
      Prob_9_0_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d[4]), Prob_9_0_sva_2, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
          {or_tmp_379 , or_tmp_380 , FOR_J_7_and_81_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_9_14_1_sva_1 <= 14'b0;
    end
    else if ( ~ FOR_J_7_or_29_rgt ) begin
      Prob_9_14_1_sva_1 <= MUX1HOT_v_14_3_2((signext_14_11(P_B_rsci_q_d[15:5])),
          Prob_9_14_1_sva_2, FOR_K_7_FOR_K_7_nor_1_psp_sva_1, {or_tmp_379 , or_tmp_380
          , FOR_J_7_and_81_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_0_sva_1_15 <= 1'b0;
    end
    else if ( ~ FOR_J_7_or_2_rgt ) begin
      Prob_0_sva_1_15 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d[15]), Prob_0_sva_2_15, (FOR_K_7_acc_7_psp_sva_1[16]),
          {or_tmp_392 , or_tmp_393 , FOR_J_7_and_27_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      FOR_J_7_and_20_cse_sva <= 1'b0;
    end
    else if ( ~ or_tmp_383 ) begin
      FOR_J_7_and_20_cse_sva <= FOR_J_7_and_stg_2_0_sva_1 & (~ (perceptron_simple_j_3_0_sva[3]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_0_sva_1_0 <= 1'b0;
    end
    else if ( ~ FOR_J_7_or_2_rgt ) begin
      Prob_0_sva_1_0 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d[4]), Prob_0_sva_2_0, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
          {or_tmp_392 , or_tmp_393 , FOR_J_7_and_27_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_0_sva_1_14_1 <= 14'b0;
    end
    else if ( ~ FOR_J_7_or_2_rgt ) begin
      Prob_0_sva_1_14_1 <= MUX1HOT_v_14_3_2((signext_14_11(P_B_rsci_q_d[15:5])),
          Prob_0_sva_2_14_1, FOR_K_7_FOR_K_7_nor_1_psp_sva_1, {or_tmp_392 , or_tmp_393
          , FOR_J_7_and_27_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_8_15_sva_1 <= 1'b0;
    end
    else if ( ~ FOR_J_7_or_26_rgt ) begin
      Prob_8_15_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d[15]), Prob_8_15_sva_2, (FOR_K_7_acc_7_psp_sva_1[16]),
          {or_tmp_405 , or_tmp_406 , FOR_J_7_and_75_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      FOR_J_7_and_19_cse_sva <= 1'b0;
    end
    else if ( ~ or_tmp_383 ) begin
      FOR_J_7_and_19_cse_sva <= FOR_J_7_and_stg_2_0_sva_1 & (perceptron_simple_j_3_0_sva[3]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_8_0_sva_1 <= 1'b0;
    end
    else if ( ~ FOR_J_7_or_26_rgt ) begin
      Prob_8_0_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d[4]), Prob_8_0_sva_2, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
          {or_tmp_405 , or_tmp_406 , FOR_J_7_and_75_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_8_14_1_sva_1 <= 14'b0;
    end
    else if ( ~ FOR_J_7_or_26_rgt ) begin
      Prob_8_14_1_sva_1 <= MUX1HOT_v_14_3_2((signext_14_11(P_B_rsci_q_d[15:5])),
          Prob_8_14_1_sva_2, FOR_K_7_FOR_K_7_nor_1_psp_sva_1, {or_tmp_405 , or_tmp_406
          , FOR_J_7_and_75_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_1_15_sva_1 <= 1'b0;
    end
    else if ( ~ FOR_J_7_or_23_rgt ) begin
      Prob_1_15_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d[15]), Prob_1_15_sva_2, (FOR_K_7_acc_7_psp_sva_1[16]),
          {or_tmp_418 , or_tmp_419 , FOR_J_7_and_69_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      FOR_J_7_and_18_cse_sva <= 1'b0;
    end
    else if ( ~ or_tmp_383 ) begin
      FOR_J_7_and_18_cse_sva <= FOR_J_7_and_stg_2_1_sva_1 & (~ (perceptron_simple_j_3_0_sva[3]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_1_0_sva_1 <= 1'b0;
    end
    else if ( ~ FOR_J_7_or_23_rgt ) begin
      Prob_1_0_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d[4]), Prob_1_0_sva_2, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
          {or_tmp_418 , or_tmp_419 , FOR_J_7_and_69_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_1_14_1_sva_1 <= 14'b0;
    end
    else if ( ~ FOR_J_7_or_23_rgt ) begin
      Prob_1_14_1_sva_1 <= MUX1HOT_v_14_3_2((signext_14_11(P_B_rsci_q_d[15:5])),
          Prob_1_14_1_sva_2, FOR_K_7_FOR_K_7_nor_1_psp_sva_1, {or_tmp_418 , or_tmp_419
          , FOR_J_7_and_69_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_7_15_sva_1 <= 1'b0;
    end
    else if ( ~ FOR_J_7_or_20_rgt ) begin
      Prob_7_15_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d[15]), Prob_7_15_sva_2, (FOR_K_7_acc_7_psp_sva_1[16]),
          {or_tmp_431 , or_tmp_432 , FOR_J_7_and_63_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      FOR_J_7_and_17_cse_sva <= 1'b0;
    end
    else if ( ~ or_tmp_383 ) begin
      FOR_J_7_and_17_cse_sva <= FOR_J_7_and_stg_1_3_sva_1 & (perceptron_simple_j_3_0_sva[3:2]==2'b01);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_7_0_sva_1 <= 1'b0;
    end
    else if ( ~ FOR_J_7_or_20_rgt ) begin
      Prob_7_0_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d[4]), Prob_7_0_sva_2, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
          {or_tmp_431 , or_tmp_432 , FOR_J_7_and_63_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_7_14_1_sva_1 <= 14'b0;
    end
    else if ( ~ FOR_J_7_or_20_rgt ) begin
      Prob_7_14_1_sva_1 <= MUX1HOT_v_14_3_2((signext_14_11(P_B_rsci_q_d[15:5])),
          Prob_7_14_1_sva_2, FOR_K_7_FOR_K_7_nor_1_psp_sva_1, {or_tmp_431 , or_tmp_432
          , FOR_J_7_and_63_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_2_15_sva_1 <= 1'b0;
    end
    else if ( ~ FOR_J_7_or_17_rgt ) begin
      Prob_2_15_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d[15]), Prob_2_15_sva_2, (FOR_K_7_acc_7_psp_sva_1[16]),
          {or_tmp_444 , or_tmp_445 , FOR_J_7_and_57_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      FOR_J_7_and_16_cse_sva <= 1'b0;
    end
    else if ( ~ or_tmp_383 ) begin
      FOR_J_7_and_16_cse_sva <= FOR_J_7_and_stg_1_2_sva_1 & (perceptron_simple_j_3_0_sva[3:2]==2'b00);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_2_0_sva_1 <= 1'b0;
    end
    else if ( ~ FOR_J_7_or_17_rgt ) begin
      Prob_2_0_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d[4]), Prob_2_0_sva_2, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
          {or_tmp_444 , or_tmp_445 , FOR_J_7_and_57_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_2_14_1_sva_1 <= 14'b0;
    end
    else if ( ~ FOR_J_7_or_17_rgt ) begin
      Prob_2_14_1_sva_1 <= MUX1HOT_v_14_3_2((signext_14_11(P_B_rsci_q_d[15:5])),
          Prob_2_14_1_sva_2, FOR_K_7_FOR_K_7_nor_1_psp_sva_1, {or_tmp_444 , or_tmp_445
          , FOR_J_7_and_57_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_6_15_sva_1 <= 1'b0;
    end
    else if ( ~ FOR_J_7_or_14_rgt ) begin
      Prob_6_15_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d[15]), Prob_6_15_sva_2, (FOR_K_7_acc_7_psp_sva_1[16]),
          {or_tmp_457 , or_tmp_458 , FOR_J_7_and_51_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      FOR_J_7_and_15_cse_sva <= 1'b0;
    end
    else if ( ~ or_tmp_383 ) begin
      FOR_J_7_and_15_cse_sva <= FOR_J_7_and_stg_1_2_sva_1 & (perceptron_simple_j_3_0_sva[3:2]==2'b01);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_6_0_sva_1 <= 1'b0;
    end
    else if ( ~ FOR_J_7_or_14_rgt ) begin
      Prob_6_0_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d[4]), Prob_6_0_sva_2, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
          {or_tmp_457 , or_tmp_458 , FOR_J_7_and_51_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_6_14_1_sva_1 <= 14'b0;
    end
    else if ( ~ FOR_J_7_or_14_rgt ) begin
      Prob_6_14_1_sva_1 <= MUX1HOT_v_14_3_2((signext_14_11(P_B_rsci_q_d[15:5])),
          Prob_6_14_1_sva_2, FOR_K_7_FOR_K_7_nor_1_psp_sva_1, {or_tmp_457 , or_tmp_458
          , FOR_J_7_and_51_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_3_15_sva_1 <= 1'b0;
    end
    else if ( ~ FOR_J_7_or_11_rgt ) begin
      Prob_3_15_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d[15]), Prob_3_15_sva_2, (FOR_K_7_acc_7_psp_sva_1[16]),
          {or_tmp_470 , or_tmp_471 , FOR_J_7_and_45_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      FOR_J_7_and_14_cse_sva <= 1'b0;
    end
    else if ( ~ or_tmp_383 ) begin
      FOR_J_7_and_14_cse_sva <= FOR_J_7_and_stg_1_3_sva_1 & (perceptron_simple_j_3_0_sva[3:2]==2'b00);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_3_0_sva_1 <= 1'b0;
    end
    else if ( ~ FOR_J_7_or_11_rgt ) begin
      Prob_3_0_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d[4]), Prob_3_0_sva_2, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
          {or_tmp_470 , or_tmp_471 , FOR_J_7_and_45_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_3_14_1_sva_1 <= 14'b0;
    end
    else if ( ~ FOR_J_7_or_11_rgt ) begin
      Prob_3_14_1_sva_1 <= MUX1HOT_v_14_3_2((signext_14_11(P_B_rsci_q_d[15:5])),
          Prob_3_14_1_sva_2, FOR_K_7_FOR_K_7_nor_1_psp_sva_1, {or_tmp_470 , or_tmp_471
          , FOR_J_7_and_45_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_5_15_sva_1 <= 1'b0;
    end
    else if ( ~ FOR_J_7_or_8_rgt ) begin
      Prob_5_15_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d[15]), Prob_5_15_sva_2, (FOR_K_7_acc_7_psp_sva_1[16]),
          {or_tmp_483 , or_tmp_484 , FOR_J_7_and_39_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      FOR_J_7_and_13_cse_sva <= 1'b0;
    end
    else if ( ~ or_tmp_383 ) begin
      FOR_J_7_and_13_cse_sva <= FOR_J_7_and_stg_1_1_sva_1 & (perceptron_simple_j_3_0_sva[3:2]==2'b01);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_5_0_sva_1 <= 1'b0;
    end
    else if ( ~ FOR_J_7_or_8_rgt ) begin
      Prob_5_0_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d[4]), Prob_5_0_sva_2, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
          {or_tmp_483 , or_tmp_484 , FOR_J_7_and_39_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_5_14_1_sva_1 <= 14'b0;
    end
    else if ( ~ FOR_J_7_or_8_rgt ) begin
      Prob_5_14_1_sva_1 <= MUX1HOT_v_14_3_2((signext_14_11(P_B_rsci_q_d[15:5])),
          Prob_5_14_1_sva_2, FOR_K_7_FOR_K_7_nor_1_psp_sva_1, {or_tmp_483 , or_tmp_484
          , FOR_J_7_and_39_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_4_15_sva_1 <= 1'b0;
    end
    else if ( ~ FOR_J_7_or_5_rgt ) begin
      Prob_4_15_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d[15]), Prob_4_15_sva_2, (FOR_K_7_acc_7_psp_sva_1[16]),
          {or_tmp_496 , or_tmp_497 , FOR_J_7_and_33_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      FOR_J_7_and_12_cse_sva <= 1'b0;
    end
    else if ( ~ or_tmp_383 ) begin
      FOR_J_7_and_12_cse_sva <= FOR_J_7_and_stg_1_0_sva_1 & (perceptron_simple_j_3_0_sva[3:2]==2'b01);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_4_0_sva_1 <= 1'b0;
    end
    else if ( ~ FOR_J_7_or_5_rgt ) begin
      Prob_4_0_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d[4]), Prob_4_0_sva_2, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
          {or_tmp_496 , or_tmp_497 , FOR_J_7_and_33_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Prob_4_14_1_sva_1 <= 14'b0;
    end
    else if ( ~ FOR_J_7_or_5_rgt ) begin
      Prob_4_14_1_sva_1 <= MUX1HOT_v_14_3_2((signext_14_11(P_B_rsci_q_d[15:5])),
          Prob_4_14_1_sva_2, FOR_K_7_FOR_K_7_nor_1_psp_sva_1, {or_tmp_496 , or_tmp_497
          , FOR_J_7_and_33_rgt});
    end
  end
  assign FOR_K_7_mux_1_nl = MUX_s_1_2_2(Prob_9_15_sva_1, (FOR_K_7_acc_7_psp_sva_1[16]),
      FOR_J_7_and_21_cse_sva);
  assign FOR_K_7_mux_2_nl = MUX_s_1_2_2(Prob_9_0_sva_1, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
      FOR_J_7_and_21_cse_sva);
  assign Prob_Prob_nor_nl = ~(FOR_J_7_and_21_cse_sva | or_tmp_125);
  assign Prob_and_19_nl = FOR_J_7_and_21_cse_sva & (~ or_tmp_125);
  assign FOR_K_7_mux_4_nl = MUX_s_1_2_2(Prob_8_15_sva_1, (FOR_K_7_acc_7_psp_sva_1[16]),
      FOR_J_7_and_19_cse_sva);
  assign FOR_K_7_mux_5_nl = MUX_s_1_2_2(Prob_8_0_sva_1, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
      FOR_J_7_and_19_cse_sva);
  assign Prob_Prob_nor_1_nl = ~(FOR_J_7_and_19_cse_sva | or_tmp_125);
  assign Prob_and_17_nl = FOR_J_7_and_19_cse_sva & (~ or_tmp_125);
  assign FOR_K_7_mux_7_nl = MUX_s_1_2_2(Prob_1_15_sva_1, (FOR_K_7_acc_7_psp_sva_1[16]),
      FOR_J_7_and_18_cse_sva);
  assign FOR_K_7_mux_8_nl = MUX_s_1_2_2(Prob_1_0_sva_1, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
      FOR_J_7_and_18_cse_sva);
  assign Prob_Prob_nor_2_nl = ~(FOR_J_7_and_18_cse_sva | or_tmp_125);
  assign Prob_and_15_nl = FOR_J_7_and_18_cse_sva & (~ or_tmp_125);
  assign FOR_K_7_mux_10_nl = MUX_s_1_2_2(Prob_7_15_sva_1, (FOR_K_7_acc_7_psp_sva_1[16]),
      FOR_J_7_and_17_cse_sva);
  assign FOR_K_7_mux_11_nl = MUX_s_1_2_2(Prob_7_0_sva_1, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
      FOR_J_7_and_17_cse_sva);
  assign Prob_Prob_nor_3_nl = ~(FOR_J_7_and_17_cse_sva | or_tmp_125);
  assign Prob_and_13_nl = FOR_J_7_and_17_cse_sva & (~ or_tmp_125);
  assign FOR_K_7_mux_13_nl = MUX_s_1_2_2(Prob_2_15_sva_1, (FOR_K_7_acc_7_psp_sva_1[16]),
      FOR_J_7_and_16_cse_sva);
  assign FOR_K_7_mux_14_nl = MUX_s_1_2_2(Prob_2_0_sva_1, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
      FOR_J_7_and_16_cse_sva);
  assign Prob_Prob_nor_4_nl = ~(FOR_J_7_and_16_cse_sva | or_tmp_125);
  assign Prob_and_11_nl = FOR_J_7_and_16_cse_sva & (~ or_tmp_125);
  assign FOR_K_7_mux_16_nl = MUX_s_1_2_2(Prob_6_15_sva_1, (FOR_K_7_acc_7_psp_sva_1[16]),
      FOR_J_7_and_15_cse_sva);
  assign FOR_K_7_mux_17_nl = MUX_s_1_2_2(Prob_6_0_sva_1, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
      FOR_J_7_and_15_cse_sva);
  assign Prob_Prob_nor_5_nl = ~(FOR_J_7_and_15_cse_sva | or_tmp_125);
  assign Prob_and_9_nl = FOR_J_7_and_15_cse_sva & (~ or_tmp_125);
  assign FOR_K_7_mux_19_nl = MUX_s_1_2_2(Prob_3_15_sva_1, (FOR_K_7_acc_7_psp_sva_1[16]),
      FOR_J_7_and_14_cse_sva);
  assign FOR_K_7_mux_20_nl = MUX_s_1_2_2(Prob_3_0_sva_1, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
      FOR_J_7_and_14_cse_sva);
  assign Prob_Prob_nor_6_nl = ~(FOR_J_7_and_14_cse_sva | or_tmp_125);
  assign Prob_and_7_nl = FOR_J_7_and_14_cse_sva & (~ or_tmp_125);
  assign FOR_K_7_mux_22_nl = MUX_s_1_2_2(Prob_5_15_sva_1, (FOR_K_7_acc_7_psp_sva_1[16]),
      FOR_J_7_and_13_cse_sva);
  assign FOR_K_7_mux_23_nl = MUX_s_1_2_2(Prob_5_0_sva_1, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
      FOR_J_7_and_13_cse_sva);
  assign Prob_Prob_nor_7_nl = ~(FOR_J_7_and_13_cse_sva | or_tmp_125);
  assign Prob_and_5_nl = FOR_J_7_and_13_cse_sva & (~ or_tmp_125);
  assign FOR_K_7_mux_25_nl = MUX_s_1_2_2(Prob_4_15_sva_1, (FOR_K_7_acc_7_psp_sva_1[16]),
      FOR_J_7_and_12_cse_sva);
  assign FOR_K_7_mux_26_nl = MUX_s_1_2_2(Prob_4_0_sva_1, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
      FOR_J_7_and_12_cse_sva);
  assign Prob_Prob_nor_8_nl = ~(FOR_J_7_and_12_cse_sva | or_tmp_125);
  assign Prob_and_3_nl = FOR_J_7_and_12_cse_sva & (~ or_tmp_125);
  assign CR1_simple_i_nor_nl = ~((fsm_output[2]) | (fsm_output[5]) | (fsm_output[6]));
  assign not_408_nl = ~ (fsm_output[27]);
  assign MP1_simple_i_N_not_nl = ~ (fsm_output[26]);
  assign MP1_simple_a_nor_nl = ~((fsm_output[25]) | (fsm_output[21]));
  assign not_404_nl = ~ (fsm_output[53]);
  assign MP2_simple_i_N_not_nl = ~ (fsm_output[52]);
  assign MP2_simple_a_nor_nl = ~((fsm_output[51]) | (fsm_output[47]));
  assign FOR_K_7_mux_28_nl = MUX_s_1_2_2(Prob_0_sva_1_15, (FOR_K_7_acc_7_psp_sva_1[16]),
      FOR_J_7_and_20_cse_sva);
  assign FOR_K_7_mux_29_nl = MUX_s_1_2_2(Prob_0_sva_1_0, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
      FOR_J_7_and_20_cse_sva);
  assign Prob_Prob_nor_9_nl = ~(FOR_J_7_and_20_cse_sva | or_tmp_376);
  assign Prob_and_1_nl = FOR_J_7_and_20_cse_sva & (~ or_tmp_376);
  assign nl_FOR_K_7_acc_nl = conv_u2s_6_7(perceptron_simple_k_7_0_sva_2[7:2]) + 7'b1010011;
  assign FOR_K_7_acc_nl = nl_FOR_K_7_acc_nl[6:0];
  assign for_mux_1_nl = MUX_s_1_2_2(max_sva_15, for_slc_Prob_16_15_0_cse_sva_15_1,
      z_out_22[16]);
  assign for_mux_2_nl = MUX_s_1_2_2(max_sva_0, for_slc_Prob_16_15_0_cse_sva_0_1,
      z_out_22[16]);
  assign CR1_simple_l_not_1_nl = ~ (fsm_output[2]);
  assign CR1_simple_j_not_nl = ~ reg_CR1_simple_l_1_6_0_sva_5_CR1_simple_l_or_cse;
  assign CR1_simple_aux_mux_14_nl = MUX_s_1_2_2(CR1_simple_aux_15_lpi_7_mx1, CR1_simple_aux_15_lpi_7_dfm,
      fsm_output[9]);
  assign CR1_simple_aux_mux_13_nl = MUX_v_14_2_2(CR1_simple_aux_14_1_lpi_7_mx1, CR1_simple_aux_14_1_lpi_7_dfm,
      fsm_output[9]);
  assign not_410_nl = ~ or_332_cse;
  assign CR1_simple_aux_mux_12_nl = MUX_s_1_2_2(CR1_simple_aux_0_lpi_7_mx1, CR1_simple_aux_0_lpi_7_dfm,
      fsm_output[9]);
  assign MP1_simple_i_not_nl = ~ (fsm_output[20]);
  assign MP1_simple_b_not_nl = ~ (fsm_output[21]);
  assign memory_1_mux_3_nl = MUX_v_16_2_2(MP1_simple_bigger_lpi_6_mx1, MP1_simple_bigger_lpi_6_dfm_1,
      fsm_output[25]);
  assign MP1_simple_bigger_not_nl = ~ (fsm_output[21]);
  assign CR1_simple_aux_mux_11_nl = MUX_s_1_2_2(CR2_simple_aux_15_lpi_7_mx1, CR2_simple_aux_15_lpi_7_dfm,
      fsm_output[35]);
  assign CR1_simple_aux_mux_10_nl = MUX_v_14_2_2(CR2_simple_aux_14_1_lpi_7_mx1, CR2_simple_aux_14_1_lpi_7_dfm,
      fsm_output[35]);
  assign not_406_nl = ~ or_400_cse;
  assign CR1_simple_aux_mux_9_nl = MUX_s_1_2_2(CR2_simple_aux_0_lpi_7_mx1, CR2_simple_aux_0_lpi_7_dfm,
      fsm_output[35]);
  assign MP2_simple_i_not_nl = ~ (fsm_output[46]);
  assign MP2_simple_b_not_nl = ~ (fsm_output[47]);
  assign memory_1_mux_4_nl = MUX_v_16_2_2(MP2_simple_bigger_lpi_6_mx1, MP2_simple_bigger_lpi_6_dfm_1,
      fsm_output[51]);
  assign MP2_simple_bigger_not_nl = ~ (fsm_output[47]);
  assign CR1_simple_aux_mux_8_nl = MUX_s_1_2_2(CR3_simple_aux_15_lpi_7_mx1, CR3_simple_aux_15_lpi_7_dfm,
      fsm_output[61]);
  assign CR1_simple_aux_mux_7_nl = MUX_v_14_2_2(CR3_simple_aux_14_1_lpi_7_mx1, CR3_simple_aux_14_1_lpi_7_dfm,
      fsm_output[61]);
  assign not_402_nl = ~ or_468_cse;
  assign CR1_simple_aux_mux_6_nl = MUX_s_1_2_2(CR3_simple_aux_0_lpi_7_mx1, CR3_simple_aux_0_lpi_7_dfm,
      fsm_output[61]);
  assign MP3_simple_i_not_nl = ~ (fsm_output[72]);
  assign MP3_simple_a_not_nl = ~ reg_MP3_simple_b_1_MP3_simple_b_or_cse;
  assign MP3_simple_b_not_nl = ~ (fsm_output[73]);
  assign memory_1_mux_5_nl = MUX_v_16_2_2(MP3_simple_bigger_lpi_6_mx1, MP3_simple_bigger_lpi_6_dfm_1,
      fsm_output[77]);
  assign MP3_simple_bigger_not_nl = ~ (fsm_output[73]);
  assign nl_reshape_simple_add_N_10_0_sva_1  = reshape_simple_add_N_10_0_lpi_4 +
      11'b1;
  assign INIT_I_or_13_nl = (fsm_output[3]) | (fsm_output[10]) | (fsm_output[15])
      | (fsm_output[5]) | (fsm_output[13]) | (fsm_output[18]);
  assign INIT_I_or_14_nl = (fsm_output[29]) | (fsm_output[36]) | (fsm_output[41])
      | (fsm_output[39]) | (fsm_output[26]) | (fsm_output[27]) | (fsm_output[31])
      | (fsm_output[44]);
  assign INIT_I_or_15_nl = (fsm_output[55]) | (fsm_output[62]) | (fsm_output[67])
      | (fsm_output[65]) | (fsm_output[52]) | (fsm_output[53]) | (fsm_output[57])
      | (fsm_output[70]);
  assign INIT_I_mux1h_7_nl = MUX1HOT_v_2_7_2((z_out_9[4:3]), (z_out_5[3:2]), (z_out_6[2:1]),
      (~ CR3_simple_a_1_0_sva), (FOR_A_1_oelse_acc_1_ncse_sva_2[3:2]), MP3_simple_i_2_1_sva,
      (FOR_A_3_oelse_acc_1_ncse_sva_2[2:1]), {(INIT_I_or_13_nl) , (INIT_I_or_14_nl)
      , (INIT_I_or_15_nl) , (fsm_output[59]) , (fsm_output[22]) , (fsm_output[74])
      , (fsm_output[48])});
  assign INIT_I_nor_1_nl = ~((fsm_output[3]) | (fsm_output[10]) | (fsm_output[15])
      | (fsm_output[29]) | (fsm_output[36]) | (fsm_output[41]) | (fsm_output[55])
      | (fsm_output[62]) | (fsm_output[67]) | (fsm_output[59]) | (fsm_output[5])
      | (fsm_output[13]) | (fsm_output[39]) | (fsm_output[65]) | (fsm_output[18])
      | (fsm_output[26]) | (fsm_output[27]) | (fsm_output[31]) | (fsm_output[44])
      | (fsm_output[52]) | (fsm_output[53]) | (fsm_output[57]) | (fsm_output[70])
      | (fsm_output[22]) | (fsm_output[48]));
  assign INIT_I_or_17_nl = (fsm_output[3]) | (fsm_output[10]) | (fsm_output[15])
      | (fsm_output[29]) | (fsm_output[36]) | (fsm_output[41]) | (fsm_output[55])
      | (fsm_output[62]) | (fsm_output[67]) | (fsm_output[5]) | (fsm_output[13])
      | (fsm_output[39]) | (fsm_output[65]) | (fsm_output[18]) | (fsm_output[26])
      | (fsm_output[27]) | (fsm_output[31]) | (fsm_output[44]) | (fsm_output[52])
      | (fsm_output[53]) | (fsm_output[57]) | (fsm_output[70]) | (fsm_output[22])
      | (fsm_output[48]);
  assign INIT_I_mux1h_8_nl = MUX1HOT_v_2_3_2(2'b1, CR3_simple_b_1_0_sva, ({1'b0 ,
      (MP3_simple_a_1_0_sva[1])}), {(INIT_I_or_17_nl) , (fsm_output[59]) , (fsm_output[74])});
  assign nl_acc_nl = ({1'b1 , (INIT_I_mux1h_7_nl) , (INIT_I_nor_1_nl)}) + conv_u2u_3_4({(INIT_I_mux1h_8_nl)
      , 1'b1});
  assign acc_nl = nl_acc_nl[3:0];
  assign z_out = readslicef_4_3_1((acc_nl));
  assign nl_FOR_A_3_if_acc_16_nl = MP2_simple_j_3_1_sva + conv_u2u_1_3(MP2_simple_b_1_0_sva[1]);
  assign FOR_A_3_if_acc_16_nl = nl_FOR_A_3_if_acc_16_nl[2:0];
  assign FOR_A_1_if_mux1h_9_nl = MUX1HOT_v_2_3_2((z_out_7[3:2]), (readslicef_3_2_1((FOR_A_3_if_acc_16_nl))),
      MP3_simple_j_2_1_sva, {(fsm_output[22]) , (fsm_output[48]) , (fsm_output[74])});
  assign FOR_A_1_if_nor_3_nl = ~((fsm_output[22]) | (fsm_output[48]));
  assign FOR_A_1_if_FOR_A_1_if_or_1_nl = (MP3_simple_b_1_0_sva[1]) | (fsm_output[22])
      | (fsm_output[48]);
  assign nl_acc_1_nl = ({1'b1 , (FOR_A_1_if_mux1h_9_nl) , (FOR_A_1_if_nor_3_nl)})
      + conv_u2u_2_4({(FOR_A_1_if_FOR_A_1_if_or_1_nl) , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[3:0];
  assign z_out_1_2 = readslicef_4_1_3((acc_1_nl));
  assign FOR_B_or_3_nl = (fsm_output[84]) | (fsm_output[81]);
  assign FOR_B_mux1h_6_nl = MUX1HOT_v_2_19_2(CR1_simple_b_1_0_sva, MP1_simple_a_1_0_sva,
      MP1_simple_b_1_0_sva, CR2_simple_b_1_0_sva, MP2_simple_a_1_0_sva, MP2_simple_b_1_0_sva,
      CR3_simple_b_1_0_sva, ({MP3_simple_j_N_1_0_sva_1_1 , MP3_simple_j_N_1_0_sva_0}),
      ({MP3_simple_i_N_1_0_sva_1_1 , MP3_simple_i_N_1_0_sva_0}), MP3_simple_a_1_0_sva,
      MP3_simple_b_1_0_sva, CR1_simple_k_1_0_sva, CR1_simple_a_1_0_sva, CR2_simple_a_1_0_sva,
      CR3_simple_a_1_0_sva, MP3_simple_j_2_1_sva, MP3_simple_i_2_1_sva, reshape_simple_i_1_0_sva,
      reshape_simple_j_1_0_sva, {(fsm_output[7]) , (fsm_output[22]) , (fsm_output[24])
      , (fsm_output[33]) , (fsm_output[48]) , (fsm_output[50]) , (fsm_output[59])
      , (fsm_output[72]) , (fsm_output[73]) , (fsm_output[74]) , (fsm_output[76])
      , (fsm_output[14]) , (fsm_output[9]) , (fsm_output[35]) , (fsm_output[61])
      , (fsm_output[79]) , (fsm_output[78]) , (fsm_output[85]) , (FOR_B_or_3_nl)});
  assign FOR_B_FOR_B_mux_1_nl = MUX_v_2_2_2(2'b1, reshape_simple_i_1_0_sva, fsm_output[81]);
  assign nl_z_out_2 = conv_u2u_2_3(FOR_B_mux1h_6_nl) + conv_u2u_2_3(FOR_B_FOR_B_mux_1_nl);
  assign z_out_2 = nl_z_out_2[2:0];
  assign FOR_B_if_or_4_nl = (fsm_output[22]) | (fsm_output[48]) | (fsm_output[74])
      | (fsm_output[76]) | (fsm_output[33]);
  assign FOR_B_if_mux1h_6_nl = MUX1HOT_v_2_3_2(CR1_simple_b_1_0_sva, (z_out_4[2:1]),
      (z_out_2[2:1]), {(fsm_output[7]) , (FOR_B_if_or_4_nl) , (fsm_output[81])});
  assign FOR_B_if_mux1h_7_nl = MUX1HOT_v_2_7_2(CR1_simple_a_1_0_sva, MP1_simple_b_1_0_sva,
      MP2_simple_b_1_0_sva, MP3_simple_b_1_0_sva, MP3_simple_j_N_1_0_sva_1, reshape_simple_i_1_0_sva,
      CR2_simple_a_1_0_sva, {(fsm_output[7]) , (fsm_output[22]) , (fsm_output[48])
      , (fsm_output[74]) , (fsm_output[76]) , (fsm_output[81]) , (fsm_output[33])});
  assign nl_z_out_3 = conv_u2u_2_3(FOR_B_if_mux1h_6_nl) + conv_u2u_2_3(FOR_B_if_mux1h_7_nl);
  assign z_out_3 = nl_z_out_3[2:0];
  assign FOR_A_1_if_mux1h_10_nl = MUX1HOT_v_2_5_2((FOR_A_1_oelse_acc_1_ncse_sva_2[3:2]),
      CR2_simple_b_1_0_sva, (FOR_A_3_oelse_acc_1_ncse_sva_2[2:1]), MP3_simple_i_2_1_sva,
      MP3_simple_i_N_1_0_sva_1, {(fsm_output[22]) , (fsm_output[33]) , (fsm_output[48])
      , (fsm_output[74]) , (fsm_output[76])});
  assign FOR_A_1_if_and_1_nl = (MP3_simple_a_1_0_sva[1]) & (~((fsm_output[22]) |
      (fsm_output[33]) | (fsm_output[48]) | (fsm_output[76])));
  assign FOR_A_1_if_mux1h_11_nl = MUX1HOT_v_2_5_2(MP1_simple_b_1_0_sva, CR2_simple_a_1_0_sva,
      MP2_simple_b_1_0_sva, MP3_simple_b_1_0_sva, MP3_simple_j_N_1_0_sva_1, {(fsm_output[22])
      , (fsm_output[33]) , (fsm_output[48]) , (fsm_output[74]) , (fsm_output[76])});
  assign nl_acc_4_nl = conv_u2u_3_4({(FOR_A_1_if_mux1h_10_nl) , (FOR_A_1_if_and_1_nl)})
      + conv_u2u_3_4({(FOR_A_1_if_mux1h_11_nl) , 1'b1});
  assign acc_4_nl = nl_acc_4_nl[3:0];
  assign z_out_4 = readslicef_4_3_1((acc_4_nl));
  assign FOR_J_1_mux1h_2_nl = MUX1HOT_v_4_12_2(MP1_simple_j_N_3_0_sva, MP1_simple_i_N_3_0_sva,
      MP1_simple_j_4_1_sva, MP1_simple_i_4_1_sva, CR2_simple_j_1_3_0_sva, CR2_simple_i_1_3_0_sva,
      CR2_simple_j_2_3_0_sva, CR2_simple_i_2_3_0_sva, CR2_simple_j_3_0_sva, CR2_simple_i_3_0_sva,
      k_sva, perceptron_simple_j_3_0_sva, {(fsm_output[20]) , (fsm_output[21]) ,
      (fsm_output[27]) , (fsm_output[26]) , (fsm_output[31]) , (fsm_output[29]) ,
      (fsm_output[39]) , (fsm_output[36]) , (fsm_output[44]) , (fsm_output[41]) ,
      (fsm_output[90]) , (fsm_output[89])});
  assign nl_z_out_5 = (FOR_J_1_mux1h_2_nl) + 4'b1;
  assign z_out_5 = nl_z_out_5[3:0];
  assign FOR_J_3_mux1h_2_nl = MUX1HOT_v_3_10_2(MP2_simple_j_N_2_0_sva, MP2_simple_i_N_2_0_sva,
      MP2_simple_j_3_1_sva, MP2_simple_i_3_1_sva, CR3_simple_j_1_2_0_sva, CR3_simple_i_1_2_0_sva,
      CR3_simple_j_2_2_0_sva, CR3_simple_i_2_2_0_sva, CR3_simple_j_2_0_sva, CR3_simple_i_2_0_sva,
      {(fsm_output[46]) , (fsm_output[47]) , (fsm_output[53]) , (fsm_output[52])
      , (fsm_output[57]) , (fsm_output[55]) , (fsm_output[65]) , (fsm_output[62])
      , (fsm_output[70]) , (fsm_output[67])});
  assign nl_z_out_6 = (FOR_J_3_mux1h_2_nl) + 3'b1;
  assign z_out_6 = nl_z_out_6[2:0];
  assign FOR_K_6_or_5_nl = (fsm_output[81]) | (fsm_output[71]) | (fsm_output[58])
      | (fsm_output[80]) | (fsm_output[90]) | (fsm_output[89]);
  assign FOR_K_6_mux1h_2_nl = MUX1HOT_v_4_6_2(4'b1011, ({1'b0 , z_out_3}), MP1_simple_j_4_1_sva,
      (CR2_simple_l_5_0_sva_4_0_1[3:0]), (CR2_simple_l_1_5_0_sva_4_0[3:0]), (MP2_simple_k_5_0_sva_4_0[3:0]),
      {(FOR_K_6_or_5_nl) , (fsm_output[7]) , (fsm_output[22]) , memory_1_or_5_cse
      , (fsm_output[29]) , (fsm_output[48])});
  assign or_nl = (fsm_output[81]) | (fsm_output[71]) | (fsm_output[58]) | (fsm_output[80]);
  assign or_663_nl = (fsm_output[29]) | (fsm_output[36]) | (fsm_output[41]) | (fsm_output[48]);
  assign mux1h_1_nl = MUX1HOT_v_3_5_2((z_out_9[4:2]), ({z_out_17 , (CR1_simple_k_1_0_sva[0])}),
      ({2'b0 , (MP1_simple_b_1_0_sva[1])}), (z_out_5[3:1]), (z_out_10[5:3]), {(or_nl)
      , (fsm_output[7]) , (fsm_output[22]) , or_tmp_376 , (or_663_nl)});
  assign nl_z_out_7 = (FOR_K_6_mux1h_2_nl) + conv_u2u_3_4(mux1h_1_nl);
  assign z_out_7 = nl_z_out_7[3:0];
  assign FOR_A_1_if_FOR_A_1_if_and_1_nl = (z_out_3[2]) & (~((fsm_output[24]) | (fsm_output[29])
      | (fsm_output[36]) | (fsm_output[41])));
  assign FOR_A_1_if_mux1h_12_nl = MUX1HOT_v_2_5_2((z_out_3[1:0]), (MP1_simple_i_N_3_0_sva_1[3:2]),
      (CR2_simple_j_1_3_0_sva[3:2]), (CR2_simple_j_2_3_0_sva[3:2]), (CR2_simple_j_3_0_sva[3:2]),
      {(fsm_output[22]) , (fsm_output[24]) , (fsm_output[29]) , (fsm_output[36])
      , (fsm_output[41])});
  assign nl_z_out_8 = FOR_A_1_if_mux1h_4_cse + conv_u2u_3_4({(FOR_A_1_if_FOR_A_1_if_and_1_nl)
      , (FOR_A_1_if_mux1h_12_nl)});
  assign z_out_8 = nl_z_out_8[3:0];
  assign INIT_J_mux1h_2_nl = MUX1HOT_v_5_10_2(CR1_simple_j_1_4_0_sva, CR1_simple_i_1_4_0_sva,
      CR1_simple_j_2_4_0_sva, CR1_simple_i_2_4_0_sva, CR1_simple_j_4_0_sva, CR1_simple_i_4_0_sva,
      CR3_simple_l_1_4_0_sva, CR3_simple_l_4_0_sva, MP3_simple_k_4_0_sva, reshape_simple_k_4_0_sva,
      {(fsm_output[5]) , (fsm_output[3]) , (fsm_output[13]) , (fsm_output[10]) ,
      (fsm_output[18]) , (fsm_output[15]) , (fsm_output[58]) , (fsm_output[71]) ,
      (fsm_output[80]) , (fsm_output[81])});
  assign nl_z_out_9 = (INIT_J_mux1h_2_nl) + 5'b1;
  assign z_out_9 = nl_z_out_9[4:0];
  assign INIT_I_or_18_nl = (fsm_output[48]) | (fsm_output[50]);
  assign INIT_I_mux1h_9_nl = MUX1HOT_v_5_7_2(CR1_simple_i_1_4_0_sva, CR1_simple_i_2_4_0_sva,
      CR1_simple_i_4_0_sva, CR2_simple_l_1_5_0_sva_4_0, CR2_simple_l_5_0_sva_4_0_1,
      MP2_simple_k_5_0_sva_4_0, CR3_simple_k_5_0_sva_4_0, {(fsm_output[3]) , (fsm_output[10])
      , (fsm_output[15]) , (fsm_output[29]) , memory_1_or_5_cse , (INIT_I_or_18_nl)
      , (fsm_output[59])});
  assign nl_FOR_A_3_if_acc_17_nl = conv_u2u_3_4(z_out_25[3:1]) + conv_u2u_3_4(MP2_simple_j_3_1_sva);
  assign FOR_A_3_if_acc_17_nl = nl_FOR_A_3_if_acc_17_nl[3:0];
  assign INIT_I_or_19_nl = (fsm_output[29]) | (fsm_output[36]) | (fsm_output[41]);
  assign INIT_I_mux1h_10_nl = MUX1HOT_v_4_5_2((z_out_12[4:1]), (z_out_23[4:1]), (FOR_A_3_if_acc_17_nl),
      z_out_26, (z_out_11[5:2]), {INIT_I_or_6_cse , (INIT_I_or_19_nl) , (fsm_output[48])
      , (fsm_output[50]) , (fsm_output[59])});
  assign nl_z_out_10 = conv_u2u_5_6(INIT_I_mux1h_9_nl) + conv_u2u_4_6(INIT_I_mux1h_10_nl);
  assign z_out_10 = nl_z_out_10[5:0];
  assign FOR_B_4_if_mux_2_nl = MUX_v_5_2_2(CR3_simple_k_5_0_sva_4_0, reshape_simple_k_4_0_sva,
      fsm_output[81]);
  assign FOR_B_4_if_mux_3_nl = MUX_v_4_2_2(({1'b0 , (CR3_simple_l_4_0_sva[4:2])}),
      ({z_out_3 , (z_out_2[0])}), fsm_output[81]);
  assign nl_z_out_11 = conv_u2u_5_6(FOR_B_4_if_mux_2_nl) + conv_u2u_4_6(FOR_B_4_if_mux_3_nl);
  assign z_out_11 = nl_z_out_11[5:0];
  assign INIT_I_mux1h_11_nl = MUX1HOT_v_5_7_2(CR1_simple_i_1_4_0_sva, CR1_simple_i_2_4_0_sva,
      CR1_simple_i_4_0_sva, CR3_simple_l_4_0_sva, MP3_simple_k_4_0_sva, CR3_simple_l_1_4_0_sva,
      reshape_simple_k_4_0_sva, {(fsm_output[3]) , (fsm_output[10]) , (fsm_output[15])
      , memory_1_or_6_cse_1 , INIT_I_or_4_cse , (fsm_output[55]) , (fsm_output[81])});
  assign INIT_I_mux1h_12_nl = MUX1HOT_v_2_7_2((CR1_simple_j_1_4_0_sva[4:3]), (CR1_simple_j_2_4_0_sva[4:3]),
      (CR1_simple_j_4_0_sva[4:3]), (z_out_20[4:3]), (z_out_21[4:3]), (INIT_I_2_acc_6_sdt_1[4:3]),
      (z_out_11[4:3]), {(fsm_output[3]) , (fsm_output[10]) , (fsm_output[15]) , memory_1_or_6_cse_1
      , INIT_I_or_4_cse , (fsm_output[55]) , (fsm_output[81])});
  assign nl_z_out_12 = (INIT_I_mux1h_11_nl) + conv_u2u_2_5(INIT_I_mux1h_12_nl);
  assign z_out_12 = nl_z_out_12[4:0];
  assign INIT_L_mux1h_2_nl = MUX1HOT_v_6_4_2(CR1_simple_l_1_6_0_sva_5_0, CR1_simple_l_6_0_sva_5_0_1,
      MP1_simple_k_6_0_sva_5_0, CR2_simple_k_6_0_sva_5_0_1, {(fsm_output[6]) , (fsm_output[19])
      , (fsm_output[28]) , (fsm_output[40])});
  assign nl_z_out_13 = conv_u2u_6_7(INIT_L_mux1h_2_nl) + 7'b1;
  assign z_out_13 = nl_z_out_13[6:0];
  assign FOR_B_mux1h_7_nl = MUX1HOT_v_2_3_2(CR1_simple_b_1_0_sva, CR2_simple_b_1_0_sva,
      CR3_simple_a_1_0_sva, {(fsm_output[7]) , (fsm_output[33]) , (fsm_output[59])});
  assign nl_z_out_14_1_0 = (FOR_B_mux1h_7_nl) + 2'b11;
  assign z_out_14_1_0 = nl_z_out_14_1_0[1:0];
  assign FOR_B_mux1h_8_nl = MUX1HOT_v_2_3_2(CR1_simple_a_1_0_sva, CR2_simple_a_1_0_sva,
      CR3_simple_b_1_0_sva, {(fsm_output[7]) , (fsm_output[33]) , (fsm_output[59])});
  assign nl_z_out_15_1_0 = (FOR_B_mux1h_8_nl) + 2'b11;
  assign z_out_15_1_0 = nl_z_out_15_1_0[1:0];
  assign FOR_B_mux1h_9_nl = MUX1HOT_v_5_6_2(CR1_simple_j_2_4_0_sva, CR2_simple_l_1_5_0_sva_4_0,
      FOR_B_2_acc_1_psp_sva_1, CR2_simple_l_5_0_sva_4_0_1, MP2_simple_k_5_0_sva_4_0,
      CR3_simple_k_5_0_sva_4_0, {(fsm_output[7]) , (fsm_output[32]) , (fsm_output[33])
      , (fsm_output[45]) , (fsm_output[54]) , (fsm_output[66])});
  assign FOR_B_or_4_nl = (fsm_output[32]) | (fsm_output[45]) | (fsm_output[54]) |
      (fsm_output[66]);
  assign FOR_B_mux1h_10_nl = MUX1HOT_v_3_3_2(({{1{z_out_14_1_0[1]}}, z_out_14_1_0}),
      3'b1, (CR2_simple_j_aux_4_0_sva_1[4:2]), {(fsm_output[7]) , (FOR_B_or_4_nl)
      , (fsm_output[33])});
  assign nl_z_out_16 = conv_u2u_5_6(FOR_B_mux1h_9_nl) + conv_s2u_3_6(FOR_B_mux1h_10_nl);
  assign z_out_16 = nl_z_out_16[5:0];
  assign FOR_B_if_mux1h_8_nl = MUX1HOT_v_2_4_2(CR1_simple_b_1_0_sva, (CR1_simple_l_6_0_sva_5_0_1[1:0]),
      (CR1_simple_l_1_6_0_sva_5_0[1:0]), (MP1_simple_k_6_0_sva_5_0[1:0]), {(fsm_output[7])
      , memory_1_or_2_cse , (fsm_output[3]) , (fsm_output[22])});
  assign FOR_B_if_mux1h_9_nl = MUX1HOT_s_1_3_2((CR1_simple_k_1_0_sva[1]), (z_out_10[5]),
      (z_out_23[4]), {(fsm_output[7]) , INIT_I_or_6_cse , (fsm_output[22])});
  assign nl_z_out_17 = (FOR_B_if_mux1h_8_nl) + conv_u2u_1_2(FOR_B_if_mux1h_9_nl);
  assign z_out_17 = nl_z_out_17[1:0];
  assign FOR_B_if_mux1h_10_nl = MUX1HOT_v_16_4_2(F_1_rsci_q_d, F_2_rsci_q_d, F_3_rsci_q_d,
      memory_1_rsci_q_d, {(fsm_output[8]) , (fsm_output[34]) , (fsm_output[60]) ,
      (fsm_output[88])});
  assign FOR_B_if_or_5_nl = (fsm_output[34]) | (fsm_output[60]);
  assign FOR_B_if_mux1h_11_nl = MUX1HOT_v_16_3_2(image_rsci_q_d, memory_2_rsci_q_d,
      P_W_rsci_q_d, {(fsm_output[8]) , (FOR_B_if_or_5_nl) , (fsm_output[88])});
  assign mul_nl = conv_u2u_32_32($signed((FOR_B_if_mux1h_10_nl)) * $signed((FOR_B_if_mux1h_11_nl)));
  assign z_out_18_31_12 = readslicef_32_20_12((mul_nl));
  assign nl_z_out_19 = ({z_out_17 , (z_out_10[4:2])}) + (CR1_simple_l_6_0_sva_5_0_1[4:0]);
  assign z_out_19 = nl_z_out_19[4:0];
  assign nl_z_out_20 = CR3_simple_l_4_0_sva + conv_u2u_4_5(z_out_26);
  assign z_out_20 = nl_z_out_20[4:0];
  assign FOR_A_5_if_mux_1_nl = MUX_v_4_2_2(z_out_25, ({z_out_3 , (z_out_4[0])}),
      fsm_output[76]);
  assign nl_z_out_21 = MP3_simple_k_4_0_sva + conv_u2u_4_5(FOR_A_5_if_mux_1_nl);
  assign z_out_21 = nl_z_out_21[4:0];
  assign FOR_I_or_3_nl = (fsm_output[11]) | (fsm_output[16]) | (fsm_output[37]) |
      (fsm_output[42]) | (fsm_output[63]) | (fsm_output[68]);
  assign FOR_I_mux1h_2_nl = MUX1HOT_v_16_6_2(memory_1_rsci_q_d, MP1_simple_bigger_lpi_6,
      MP2_simple_bigger_lpi_6, ({1'b1 , (signext_15_3(~ (CR3_simple_j_aux_3_0_sva_1[3:1])))}),
      MP3_simple_bigger_lpi_6, ({max_sva_15 , max_sva_14_1 , max_sva_0}), {(FOR_I_or_3_nl)
      , (fsm_output[23]) , (fsm_output[49]) , (fsm_output[59]) , (fsm_output[75])
      , (fsm_output[90])});
  assign FOR_I_nor_5_nl = ~((fsm_output[11]) | (fsm_output[16]) | (fsm_output[37])
      | (fsm_output[42]) | (fsm_output[59]) | (fsm_output[63]) | (fsm_output[68]));
  assign FOR_I_or_5_nl = (fsm_output[23]) | (fsm_output[49]) | (fsm_output[75]);
  assign FOR_I_mux1h_3_nl = MUX1HOT_v_16_9_2(({CR1_simple_aux_15_lpi_7_dfm , CR1_simple_aux_14_1_lpi_7_dfm
      , CR1_simple_aux_0_lpi_7_dfm}), ({{1{BIAS_I_slc_15_1_itm[14]}}, BIAS_I_slc_15_1_itm}),
      (~ memory_1_rsci_q_d), ({CR2_simple_aux_15_lpi_7_dfm , CR2_simple_aux_14_1_lpi_7_dfm
      , CR2_simple_aux_0_lpi_7_dfm}), ({{1{BIAS_I_1_slc_15_1_itm[14]}}, BIAS_I_1_slc_15_1_itm}),
      16'b11, ({CR3_simple_aux_15_lpi_7_dfm , CR3_simple_aux_14_1_lpi_7_dfm , CR3_simple_aux_0_lpi_7_dfm}),
      ({{1{BIAS_I_2_slc_15_1_itm[14]}}, BIAS_I_2_slc_15_1_itm}), ({(~ for_slc_Prob_16_15_0_cse_sva_15_1)
      , (~ for_slc_Prob_16_15_0_cse_sva_14_1_1) , (~ for_slc_Prob_16_15_0_cse_sva_0_1)}),
      {(fsm_output[11]) , (fsm_output[16]) , (FOR_I_or_5_nl) , (fsm_output[37]) ,
      (fsm_output[42]) , (fsm_output[59]) , (fsm_output[63]) , (fsm_output[68]) ,
      (fsm_output[90])});
  assign nl_acc_21_nl = conv_s2u_17_18({(FOR_I_mux1h_2_nl) , (FOR_I_nor_5_nl)}) +
      conv_s2u_17_18({(FOR_I_mux1h_3_nl) , 1'b1});
  assign acc_21_nl = nl_acc_21_nl[17:0];
  assign z_out_22 = readslicef_18_17_1((acc_21_nl));
  assign nl_z_out_23 = conv_u2u_4_5(FOR_A_1_if_mux1h_4_cse) + conv_u2u_3_5(z_out_8[3:1]);
  assign z_out_23 = nl_z_out_23[4:0];
  assign FOR_B_2_if_mux_4_nl = MUX_s_1_2_2(CR2_simple_aux_15_lpi_7, CR3_simple_aux_15_lpi_7,
      fsm_output[60]);
  assign FOR_B_2_if_mux_5_nl = MUX_v_14_2_2(CR2_simple_aux_14_1_lpi_7, CR3_simple_aux_14_1_lpi_7,
      fsm_output[60]);
  assign FOR_B_2_if_mux_6_nl = MUX_s_1_2_2(CR2_simple_aux_0_lpi_7, CR3_simple_aux_0_lpi_7,
      fsm_output[60]);
  assign nl_z_out_24 = z_out_18_31_12 + conv_s2u_16_20({(FOR_B_2_if_mux_4_nl) , (FOR_B_2_if_mux_5_nl)
      , (FOR_B_2_if_mux_6_nl)});
  assign z_out_24 = nl_z_out_24[19:0];
  assign nl_FOR_A_5_if_acc_21_nl = MP3_simple_j_2_1_sva + conv_u2u_1_2(MP3_simple_j_2_1_sva[1]);
  assign FOR_A_5_if_acc_21_nl = nl_FOR_A_5_if_acc_21_nl[1:0];
  assign FOR_A_3_if_mux_2_nl = MUX_v_3_2_2(z_out_3, ({(FOR_A_5_if_acc_21_nl) , (MP3_simple_j_2_1_sva[0])}),
      fsm_output[74]);
  assign FOR_A_3_if_mux_3_nl = MUX_v_3_2_2(MP2_simple_j_3_1_sva, z_out_3, fsm_output[74]);
  assign nl_z_out_25 = conv_u2u_3_4(FOR_A_3_if_mux_2_nl) + conv_u2u_3_4(FOR_A_3_if_mux_3_nl);
  assign z_out_25 = nl_z_out_25[3:0];
  assign FOR_B_3_if_mux1h_2_nl = MUX1HOT_v_3_4_2(MP2_simple_j_N_2_0_sva_1, CR3_simple_i_1_2_0_sva,
      CR3_simple_i_2_2_0_sva, CR3_simple_i_2_0_sva, {(fsm_output[50]) , (fsm_output[55])
      , (fsm_output[62]) , (fsm_output[67])});
  assign FOR_B_3_if_or_1_nl = (fsm_output[55]) | (fsm_output[62]) | (fsm_output[67]);
  assign FOR_B_3_if_FOR_B_3_if_mux_1_nl = MUX_v_2_2_2((FOR_B_3_if_acc_sdt_1[2:1]),
      (z_out_27_2_0[2:1]), FOR_B_3_if_or_1_nl);
  assign nl_z_out_26 = conv_u2u_3_4(FOR_B_3_if_mux1h_2_nl) + conv_u2u_2_4(FOR_B_3_if_FOR_B_3_if_mux_1_nl);
  assign z_out_26 = nl_z_out_26[3:0];
  assign INIT_I_2_mux1h_2_nl = MUX1HOT_v_3_3_2(CR3_simple_i_1_2_0_sva, CR3_simple_i_2_2_0_sva,
      CR3_simple_i_2_0_sva, {(fsm_output[55]) , (fsm_output[62]) , (fsm_output[67])});
  assign INIT_I_2_mux1h_3_nl = MUX1HOT_v_2_3_2((CR3_simple_j_1_2_0_sva[2:1]), (CR3_simple_j_2_2_0_sva[2:1]),
      (CR3_simple_j_2_0_sva[2:1]), {(fsm_output[55]) , (fsm_output[62]) , (fsm_output[67])});
  assign nl_z_out_27_2_0 = (INIT_I_2_mux1h_2_nl) + conv_u2u_2_3(INIT_I_2_mux1h_3_nl);
  assign z_out_27_2_0 = nl_z_out_27_2_0[2:0];

  function automatic [0:0] MUX1HOT_s_1_10_2;
    input [0:0] input_9;
    input [0:0] input_8;
    input [0:0] input_7;
    input [0:0] input_6;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [9:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    result = result | ( input_6 & {1{sel[6]}});
    result = result | ( input_7 & {1{sel[7]}});
    result = result | ( input_8 & {1{sel[8]}});
    result = result | ( input_9 & {1{sel[9]}});
    MUX1HOT_s_1_10_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_5_2;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [4:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_7_2;
    input [0:0] input_6;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [6:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    result = result | ( input_6 & {1{sel[6]}});
    MUX1HOT_s_1_7_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_8_2;
    input [0:0] input_7;
    input [0:0] input_6;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [7:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    result = result | ( input_6 & {1{sel[6]}});
    result = result | ( input_7 & {1{sel[7]}});
    MUX1HOT_s_1_8_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_9_2;
    input [0:0] input_8;
    input [0:0] input_7;
    input [0:0] input_6;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [8:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    result = result | ( input_6 & {1{sel[6]}});
    result = result | ( input_7 & {1{sel[7]}});
    result = result | ( input_8 & {1{sel[8]}});
    MUX1HOT_s_1_9_2 = result;
  end
  endfunction


  function automatic [13:0] MUX1HOT_v_14_3_2;
    input [13:0] input_2;
    input [13:0] input_1;
    input [13:0] input_0;
    input [2:0] sel;
    reg [13:0] result;
  begin
    result = input_0 & {14{sel[0]}};
    result = result | ( input_1 & {14{sel[1]}});
    result = result | ( input_2 & {14{sel[2]}});
    MUX1HOT_v_14_3_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_3_2;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [2:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    MUX1HOT_v_16_3_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_4_2;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [3:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    result = result | ( input_3 & {16{sel[3]}});
    MUX1HOT_v_16_4_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_6_2;
    input [15:0] input_5;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [5:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    result = result | ( input_3 & {16{sel[3]}});
    result = result | ( input_4 & {16{sel[4]}});
    result = result | ( input_5 & {16{sel[5]}});
    MUX1HOT_v_16_6_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_9_2;
    input [15:0] input_8;
    input [15:0] input_7;
    input [15:0] input_6;
    input [15:0] input_5;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [8:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    result = result | ( input_3 & {16{sel[3]}});
    result = result | ( input_4 & {16{sel[4]}});
    result = result | ( input_5 & {16{sel[5]}});
    result = result | ( input_6 & {16{sel[6]}});
    result = result | ( input_7 & {16{sel[7]}});
    result = result | ( input_8 & {16{sel[8]}});
    MUX1HOT_v_16_9_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_19_2;
    input [1:0] input_18;
    input [1:0] input_17;
    input [1:0] input_16;
    input [1:0] input_15;
    input [1:0] input_14;
    input [1:0] input_13;
    input [1:0] input_12;
    input [1:0] input_11;
    input [1:0] input_10;
    input [1:0] input_9;
    input [1:0] input_8;
    input [1:0] input_7;
    input [1:0] input_6;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [18:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    result = result | ( input_3 & {2{sel[3]}});
    result = result | ( input_4 & {2{sel[4]}});
    result = result | ( input_5 & {2{sel[5]}});
    result = result | ( input_6 & {2{sel[6]}});
    result = result | ( input_7 & {2{sel[7]}});
    result = result | ( input_8 & {2{sel[8]}});
    result = result | ( input_9 & {2{sel[9]}});
    result = result | ( input_10 & {2{sel[10]}});
    result = result | ( input_11 & {2{sel[11]}});
    result = result | ( input_12 & {2{sel[12]}});
    result = result | ( input_13 & {2{sel[13]}});
    result = result | ( input_14 & {2{sel[14]}});
    result = result | ( input_15 & {2{sel[15]}});
    result = result | ( input_16 & {2{sel[16]}});
    result = result | ( input_17 & {2{sel[17]}});
    result = result | ( input_18 & {2{sel[18]}});
    MUX1HOT_v_2_19_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_4_2;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [3:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    result = result | ( input_3 & {2{sel[3]}});
    MUX1HOT_v_2_4_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_5_2;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [4:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    result = result | ( input_3 & {2{sel[3]}});
    result = result | ( input_4 & {2{sel[4]}});
    MUX1HOT_v_2_5_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_7_2;
    input [1:0] input_6;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [6:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    result = result | ( input_3 & {2{sel[3]}});
    result = result | ( input_4 & {2{sel[4]}});
    result = result | ( input_5 & {2{sel[5]}});
    result = result | ( input_6 & {2{sel[6]}});
    MUX1HOT_v_2_7_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_10_2;
    input [2:0] input_9;
    input [2:0] input_8;
    input [2:0] input_7;
    input [2:0] input_6;
    input [2:0] input_5;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [9:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    result = result | ( input_3 & {3{sel[3]}});
    result = result | ( input_4 & {3{sel[4]}});
    result = result | ( input_5 & {3{sel[5]}});
    result = result | ( input_6 & {3{sel[6]}});
    result = result | ( input_7 & {3{sel[7]}});
    result = result | ( input_8 & {3{sel[8]}});
    result = result | ( input_9 & {3{sel[9]}});
    MUX1HOT_v_3_10_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_4_2;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [3:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    result = result | ( input_3 & {3{sel[3]}});
    MUX1HOT_v_3_4_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_5_2;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [4:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    result = result | ( input_3 & {3{sel[3]}});
    result = result | ( input_4 & {3{sel[4]}});
    MUX1HOT_v_3_5_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_12_2;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [11:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    result = result | ( input_4 & {4{sel[4]}});
    result = result | ( input_5 & {4{sel[5]}});
    result = result | ( input_6 & {4{sel[6]}});
    result = result | ( input_7 & {4{sel[7]}});
    result = result | ( input_8 & {4{sel[8]}});
    result = result | ( input_9 & {4{sel[9]}});
    result = result | ( input_10 & {4{sel[10]}});
    result = result | ( input_11 & {4{sel[11]}});
    MUX1HOT_v_4_12_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_5_2;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [4:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    result = result | ( input_4 & {4{sel[4]}});
    MUX1HOT_v_4_5_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_6_2;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [5:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    result = result | ( input_4 & {4{sel[4]}});
    result = result | ( input_5 & {4{sel[5]}});
    MUX1HOT_v_4_6_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_7_2;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [6:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    result = result | ( input_4 & {4{sel[4]}});
    result = result | ( input_5 & {4{sel[5]}});
    result = result | ( input_6 & {4{sel[6]}});
    MUX1HOT_v_4_7_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_10_2;
    input [4:0] input_9;
    input [4:0] input_8;
    input [4:0] input_7;
    input [4:0] input_6;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [9:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | ( input_1 & {5{sel[1]}});
    result = result | ( input_2 & {5{sel[2]}});
    result = result | ( input_3 & {5{sel[3]}});
    result = result | ( input_4 & {5{sel[4]}});
    result = result | ( input_5 & {5{sel[5]}});
    result = result | ( input_6 & {5{sel[6]}});
    result = result | ( input_7 & {5{sel[7]}});
    result = result | ( input_8 & {5{sel[8]}});
    result = result | ( input_9 & {5{sel[9]}});
    MUX1HOT_v_5_10_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_6_2;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [5:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | ( input_1 & {5{sel[1]}});
    result = result | ( input_2 & {5{sel[2]}});
    result = result | ( input_3 & {5{sel[3]}});
    result = result | ( input_4 & {5{sel[4]}});
    result = result | ( input_5 & {5{sel[5]}});
    MUX1HOT_v_5_6_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_7_2;
    input [4:0] input_6;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [6:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | ( input_1 & {5{sel[1]}});
    result = result | ( input_2 & {5{sel[2]}});
    result = result | ( input_3 & {5{sel[3]}});
    result = result | ( input_4 & {5{sel[4]}});
    result = result | ( input_5 & {5{sel[5]}});
    result = result | ( input_6 & {5{sel[6]}});
    MUX1HOT_v_5_7_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_4_2;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [3:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    result = result | ( input_3 & {6{sel[3]}});
    MUX1HOT_v_6_4_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_10_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] input_2;
    input [0:0] input_3;
    input [0:0] input_4;
    input [0:0] input_5;
    input [0:0] input_6;
    input [0:0] input_7;
    input [0:0] input_8;
    input [0:0] input_9;
    input [3:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      default : begin
        result = input_9;
      end
    endcase
    MUX_s_1_10_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_10_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input [13:0] input_2;
    input [13:0] input_3;
    input [13:0] input_4;
    input [13:0] input_5;
    input [13:0] input_6;
    input [13:0] input_7;
    input [13:0] input_8;
    input [13:0] input_9;
    input [3:0] sel;
    reg [13:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      default : begin
        result = input_9;
      end
    endcase
    MUX_v_14_10_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_2_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input [0:0] sel;
    reg [13:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_14_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_14_1_13;
    input [13:0] vector;
    reg [13:0] tmp;
  begin
    tmp = vector >> 13;
    readslicef_14_1_13 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_15_1_14;
    input [14:0] vector;
    reg [14:0] tmp;
  begin
    tmp = vector >> 14;
    readslicef_15_1_14 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_16_1_15;
    input [15:0] vector;
    reg [15:0] tmp;
  begin
    tmp = vector >> 15;
    readslicef_16_1_15 = tmp[0:0];
  end
  endfunction


  function automatic [16:0] readslicef_18_17_1;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_18_17_1 = tmp[16:0];
  end
  endfunction


  function automatic [19:0] readslicef_32_20_12;
    input [31:0] vector;
    reg [31:0] tmp;
  begin
    tmp = vector >> 12;
    readslicef_32_20_12 = tmp[19:0];
  end
  endfunction


  function automatic [1:0] readslicef_3_2_1;
    input [2:0] vector;
    reg [2:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_3_2_1 = tmp[1:0];
  end
  endfunction


  function automatic [0:0] readslicef_4_1_3;
    input [3:0] vector;
    reg [3:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_4_1_3 = tmp[0:0];
  end
  endfunction


  function automatic [2:0] readslicef_4_3_1;
    input [3:0] vector;
    reg [3:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_4_3_1 = tmp[2:0];
  end
  endfunction


  function automatic [0:0] readslicef_7_1_6;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_7_1_6 = tmp[0:0];
  end
  endfunction


  function automatic [12:0] signext_13_3;
    input [2:0] vector;
  begin
    signext_13_3= {{10{vector[2]}}, vector};
  end
  endfunction


  function automatic [13:0] signext_14_1;
    input [0:0] vector;
  begin
    signext_14_1= {{13{vector[0]}}, vector};
  end
  endfunction


  function automatic [13:0] signext_14_11;
    input [10:0] vector;
  begin
    signext_14_11= {{3{vector[10]}}, vector};
  end
  endfunction


  function automatic [13:0] signext_14_3;
    input [2:0] vector;
  begin
    signext_14_3= {{11{vector[2]}}, vector};
  end
  endfunction


  function automatic [14:0] signext_15_3;
    input [2:0] vector;
  begin
    signext_15_3= {{12{vector[2]}}, vector};
  end
  endfunction


  function automatic [3:0] conv_s2s_2_4 ;
    input [1:0]  vector ;
  begin
    conv_s2s_2_4 = {{2{vector[1]}}, vector};
  end
  endfunction


  function automatic [4:0] conv_s2s_2_5 ;
    input [1:0]  vector ;
  begin
    conv_s2s_2_5 = {{3{vector[1]}}, vector};
  end
  endfunction


  function automatic [5:0] conv_s2s_2_6 ;
    input [1:0]  vector ;
  begin
    conv_s2s_2_6 = {{4{vector[1]}}, vector};
  end
  endfunction


  function automatic [3:0] conv_s2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_s2s_3_4 = {vector[2], vector};
  end
  endfunction


  function automatic [4:0] conv_s2s_3_5 ;
    input [2:0]  vector ;
  begin
    conv_s2s_3_5 = {{2{vector[2]}}, vector};
  end
  endfunction


  function automatic [5:0] conv_s2s_3_6 ;
    input [2:0]  vector ;
  begin
    conv_s2s_3_6 = {{3{vector[2]}}, vector};
  end
  endfunction


  function automatic [4:0] conv_s2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_s2s_4_5 = {vector[3], vector};
  end
  endfunction


  function automatic [6:0] conv_s2s_5_7 ;
    input [4:0]  vector ;
  begin
    conv_s2s_5_7 = {{2{vector[4]}}, vector};
  end
  endfunction


  function automatic [3:0] conv_s2u_2_4 ;
    input [1:0]  vector ;
  begin
    conv_s2u_2_4 = {{2{vector[1]}}, vector};
  end
  endfunction


  function automatic [4:0] conv_s2u_2_5 ;
    input [1:0]  vector ;
  begin
    conv_s2u_2_5 = {{3{vector[1]}}, vector};
  end
  endfunction


  function automatic [5:0] conv_s2u_3_6 ;
    input [2:0]  vector ;
  begin
    conv_s2u_3_6 = {{3{vector[2]}}, vector};
  end
  endfunction


  function automatic [4:0] conv_s2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_s2u_4_5 = {vector[3], vector};
  end
  endfunction


  function automatic [5:0] conv_s2u_4_6 ;
    input [3:0]  vector ;
  begin
    conv_s2u_4_6 = {{2{vector[3]}}, vector};
  end
  endfunction


  function automatic [5:0] conv_s2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_s2u_5_6 = {vector[4], vector};
  end
  endfunction


  function automatic [6:0] conv_s2u_5_7 ;
    input [4:0]  vector ;
  begin
    conv_s2u_5_7 = {{2{vector[4]}}, vector};
  end
  endfunction


  function automatic [6:0] conv_s2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_s2u_6_7 = {vector[5], vector};
  end
  endfunction


  function automatic [16:0] conv_s2u_16_17 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_17 = {vector[15], vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_16_19 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_19 = {{3{vector[15]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2u_16_20 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_20 = {{4{vector[15]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_17_18 ;
    input [16:0]  vector ;
  begin
    conv_s2u_17_18 = {vector[16], vector};
  end
  endfunction


  function automatic [3:0] conv_u2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2s_3_4 =  {1'b0, vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function automatic [5:0] conv_u2s_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2s_5_6 =  {1'b0, vector};
  end
  endfunction


  function automatic [6:0] conv_u2s_5_7 ;
    input [4:0]  vector ;
  begin
    conv_u2s_5_7 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [6:0] conv_u2s_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2s_6_7 =  {1'b0, vector};
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction


  function automatic [2:0] conv_u2u_1_3 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_3 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_1_4 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_4 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_2_4 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_4 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_2_5 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_5 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_3_5 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_5 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [5:0] conv_u2u_3_6 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_6 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_3_8 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_8 = {{5{1'b0}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function automatic [5:0] conv_u2u_4_6 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_6 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_4_7 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_7 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [5:0] conv_u2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_6 = {1'b0, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_6_8 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_8 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [31:0] conv_u2u_32_32 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_32 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    CNN_main_simple
// ------------------------------------------------------------------


module CNN_main_simple (
  clk, rst, image_rsc_radr, image_rsc_q, image_rsc_re, image_rsc_triosy_lz, F_1_rsc_radr,
      F_1_rsc_q, F_1_rsc_re, F_1_rsc_triosy_lz, B_1_rsc_radr, B_1_rsc_q, B_1_rsc_re,
      B_1_rsc_triosy_lz, F_2_rsc_radr, F_2_rsc_q, F_2_rsc_re, F_2_rsc_triosy_lz,
      B_2_rsc_radr, B_2_rsc_q, B_2_rsc_re, B_2_rsc_triosy_lz, F_3_rsc_radr, F_3_rsc_q,
      F_3_rsc_re, F_3_rsc_triosy_lz, B_3_rsc_radr, B_3_rsc_q, B_3_rsc_re, B_3_rsc_triosy_lz,
      P_W_rsc_radr, P_W_rsc_q, P_W_rsc_re, P_W_rsc_triosy_lz, P_B_rsc_radr, P_B_rsc_q,
      P_B_rsc_re, P_B_rsc_triosy_lz, index_rsc_dat, index_rsc_triosy_lz
);
  input clk;
  input rst;
  output [10:0] image_rsc_radr;
  input [15:0] image_rsc_q;
  output image_rsc_re;
  output image_rsc_triosy_lz;
  output [10:0] F_1_rsc_radr;
  input [15:0] F_1_rsc_q;
  output F_1_rsc_re;
  output F_1_rsc_triosy_lz;
  output [5:0] B_1_rsc_radr;
  input [15:0] B_1_rsc_q;
  output B_1_rsc_re;
  output B_1_rsc_triosy_lz;
  output [14:0] F_2_rsc_radr;
  input [15:0] F_2_rsc_q;
  output F_2_rsc_re;
  output F_2_rsc_triosy_lz;
  output [4:0] B_2_rsc_radr;
  input [15:0] B_2_rsc_q;
  output B_2_rsc_re;
  output B_2_rsc_triosy_lz;
  output [12:0] F_3_rsc_radr;
  input [15:0] F_3_rsc_q;
  output F_3_rsc_re;
  output F_3_rsc_triosy_lz;
  output [4:0] B_3_rsc_radr;
  input [15:0] B_3_rsc_q;
  output B_3_rsc_re;
  output B_3_rsc_triosy_lz;
  output [10:0] P_W_rsc_radr;
  input [15:0] P_W_rsc_q;
  output P_W_rsc_re;
  output P_W_rsc_triosy_lz;
  output [3:0] P_B_rsc_radr;
  input [15:0] P_B_rsc_q;
  output P_B_rsc_re;
  output P_B_rsc_triosy_lz;
  output [3:0] index_rsc_dat;
  output index_rsc_triosy_lz;


  // Interconnect Declarations
  wire [10:0] image_rsci_radr_d;
  wire [15:0] image_rsci_q_d;
  wire [10:0] F_1_rsci_radr_d;
  wire [15:0] F_1_rsci_q_d;
  wire [5:0] B_1_rsci_radr_d;
  wire B_1_rsci_re_d;
  wire [15:0] B_1_rsci_q_d;
  wire [14:0] F_2_rsci_radr_d;
  wire F_2_rsci_re_d;
  wire [15:0] F_2_rsci_q_d;
  wire [4:0] B_2_rsci_radr_d;
  wire B_2_rsci_re_d;
  wire [15:0] B_2_rsci_q_d;
  wire [12:0] F_3_rsci_radr_d;
  wire F_3_rsci_re_d;
  wire [15:0] F_3_rsci_q_d;
  wire [4:0] B_3_rsci_radr_d;
  wire B_3_rsci_re_d;
  wire [15:0] B_3_rsci_q_d;
  wire [10:0] P_W_rsci_radr_d;
  wire P_W_rsci_re_d;
  wire [15:0] P_W_rsci_q_d;
  wire [3:0] P_B_rsci_radr_d;
  wire P_B_rsci_re_d;
  wire [15:0] P_B_rsci_q_d;
  wire [10:0] memory_1_rsci_radr_d;
  wire [10:0] memory_1_rsci_wadr_d;
  wire [15:0] memory_1_rsci_d_d;
  wire memory_1_rsci_we_d;
  wire memory_1_rsci_re_d;
  wire [15:0] memory_1_rsci_q_d;
  wire [10:0] memory_2_rsci_radr_d;
  wire [10:0] memory_2_rsci_wadr_d;
  wire [15:0] memory_2_rsci_d_d;
  wire memory_2_rsci_we_d;
  wire memory_2_rsci_re_d;
  wire [15:0] memory_2_rsci_q_d;
  wire memory_1_rsc_we;
  wire [15:0] memory_1_rsc_d;
  wire [10:0] memory_1_rsc_wadr;
  wire memory_1_rsc_re;
  wire [15:0] memory_1_rsc_q;
  wire [10:0] memory_1_rsc_radr;
  wire memory_2_rsc_we;
  wire [15:0] memory_2_rsc_d;
  wire [10:0] memory_2_rsc_wadr;
  wire memory_2_rsc_re;
  wire [15:0] memory_2_rsc_q;
  wire [10:0] memory_2_rsc_radr;
  wire image_rsci_re_d_iff;


  // Interconnect Declarations for Component Instantiations 
  BLOCK_1R1W_RBW #(.data_width(32'sd16),
  .addr_width(32'sd11),
  .depth(32'sd1728)) memory_1_rsc_comp (
      .radr(memory_1_rsc_radr),
      .wadr(memory_1_rsc_wadr),
      .d(memory_1_rsc_d),
      .we(memory_1_rsc_we),
      .re(memory_1_rsc_re),
      .clk(clk),
      .q(memory_1_rsc_q)
    );
  BLOCK_1R1W_RBW #(.data_width(32'sd16),
  .addr_width(32'sd11),
  .depth(32'sd1728)) memory_2_rsc_comp (
      .radr(memory_2_rsc_radr),
      .wadr(memory_2_rsc_wadr),
      .d(memory_2_rsc_d),
      .we(memory_2_rsc_we),
      .re(memory_2_rsc_re),
      .clk(clk),
      .q(memory_2_rsc_q)
    );
  CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1728_1_gen image_rsci (
      .re(image_rsc_re),
      .q(image_rsc_q),
      .radr(image_rsc_radr),
      .radr_d(image_rsci_radr_d),
      .re_d(image_rsci_re_d_iff),
      .q_d(image_rsci_q_d)
    );
  CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1728_2_gen F_1_rsci (
      .re(F_1_rsc_re),
      .q(F_1_rsc_q),
      .radr(F_1_rsc_radr),
      .radr_d(F_1_rsci_radr_d),
      .re_d(image_rsci_re_d_iff),
      .q_d(F_1_rsci_q_d)
    );
  CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_6_64_3_gen B_1_rsci (
      .re(B_1_rsc_re),
      .q(B_1_rsc_q),
      .radr(B_1_rsc_radr),
      .radr_d(B_1_rsci_radr_d),
      .re_d(B_1_rsci_re_d),
      .q_d(B_1_rsci_q_d)
    );
  CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_15_18432_4_gen F_2_rsci (
      .re(F_2_rsc_re),
      .q(F_2_rsc_q),
      .radr(F_2_rsc_radr),
      .radr_d(F_2_rsci_radr_d),
      .re_d(F_2_rsci_re_d),
      .q_d(F_2_rsci_q_d)
    );
  CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_5_32_5_gen B_2_rsci (
      .re(B_2_rsc_re),
      .q(B_2_rsc_q),
      .radr(B_2_rsc_radr),
      .radr_d(B_2_rsci_radr_d),
      .re_d(B_2_rsci_re_d),
      .q_d(B_2_rsci_q_d)
    );
  CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_13_5760_6_gen F_3_rsci (
      .re(F_3_rsc_re),
      .q(F_3_rsc_q),
      .radr(F_3_rsc_radr),
      .radr_d(F_3_rsci_radr_d),
      .re_d(F_3_rsci_re_d),
      .q_d(F_3_rsci_q_d)
    );
  CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_5_20_7_gen B_3_rsci (
      .re(B_3_rsc_re),
      .q(B_3_rsc_q),
      .radr(B_3_rsc_radr),
      .radr_d(B_3_rsci_radr_d),
      .re_d(B_3_rsci_re_d),
      .q_d(B_3_rsci_q_d)
    );
  CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1800_8_gen P_W_rsci (
      .re(P_W_rsc_re),
      .q(P_W_rsc_q),
      .radr(P_W_rsc_radr),
      .radr_d(P_W_rsci_radr_d),
      .re_d(P_W_rsci_re_d),
      .q_d(P_W_rsci_q_d)
    );
  CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_4_10_9_gen P_B_rsci (
      .re(P_B_rsc_re),
      .q(P_B_rsc_q),
      .radr(P_B_rsc_radr),
      .radr_d(P_B_rsci_radr_d),
      .re_d(P_B_rsci_re_d),
      .q_d(P_B_rsci_q_d)
    );
  CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_11_1728_11_gen memory_1_rsci
      (
      .we(memory_1_rsc_we),
      .d(memory_1_rsc_d),
      .wadr(memory_1_rsc_wadr),
      .re(memory_1_rsc_re),
      .q(memory_1_rsc_q),
      .radr(memory_1_rsc_radr),
      .radr_d(memory_1_rsci_radr_d),
      .wadr_d(memory_1_rsci_wadr_d),
      .d_d(memory_1_rsci_d_d),
      .we_d(memory_1_rsci_we_d),
      .re_d(memory_1_rsci_re_d),
      .q_d(memory_1_rsci_q_d)
    );
  CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_11_1728_12_gen memory_2_rsci
      (
      .we(memory_2_rsc_we),
      .d(memory_2_rsc_d),
      .wadr(memory_2_rsc_wadr),
      .re(memory_2_rsc_re),
      .q(memory_2_rsc_q),
      .radr(memory_2_rsc_radr),
      .radr_d(memory_2_rsci_radr_d),
      .wadr_d(memory_2_rsci_wadr_d),
      .d_d(memory_2_rsci_d_d),
      .we_d(memory_2_rsci_we_d),
      .re_d(memory_2_rsci_re_d),
      .q_d(memory_2_rsci_q_d)
    );
  CNN_main_simple_core CNN_main_simple_core_inst (
      .clk(clk),
      .rst(rst),
      .image_rsc_triosy_lz(image_rsc_triosy_lz),
      .F_1_rsc_triosy_lz(F_1_rsc_triosy_lz),
      .B_1_rsc_triosy_lz(B_1_rsc_triosy_lz),
      .F_2_rsc_triosy_lz(F_2_rsc_triosy_lz),
      .B_2_rsc_triosy_lz(B_2_rsc_triosy_lz),
      .F_3_rsc_triosy_lz(F_3_rsc_triosy_lz),
      .B_3_rsc_triosy_lz(B_3_rsc_triosy_lz),
      .P_W_rsc_triosy_lz(P_W_rsc_triosy_lz),
      .P_B_rsc_triosy_lz(P_B_rsc_triosy_lz),
      .index_rsc_dat(index_rsc_dat),
      .index_rsc_triosy_lz(index_rsc_triosy_lz),
      .image_rsci_radr_d(image_rsci_radr_d),
      .image_rsci_q_d(image_rsci_q_d),
      .F_1_rsci_radr_d(F_1_rsci_radr_d),
      .F_1_rsci_q_d(F_1_rsci_q_d),
      .B_1_rsci_radr_d(B_1_rsci_radr_d),
      .B_1_rsci_re_d(B_1_rsci_re_d),
      .B_1_rsci_q_d(B_1_rsci_q_d),
      .F_2_rsci_radr_d(F_2_rsci_radr_d),
      .F_2_rsci_re_d(F_2_rsci_re_d),
      .F_2_rsci_q_d(F_2_rsci_q_d),
      .B_2_rsci_radr_d(B_2_rsci_radr_d),
      .B_2_rsci_re_d(B_2_rsci_re_d),
      .B_2_rsci_q_d(B_2_rsci_q_d),
      .F_3_rsci_radr_d(F_3_rsci_radr_d),
      .F_3_rsci_re_d(F_3_rsci_re_d),
      .F_3_rsci_q_d(F_3_rsci_q_d),
      .B_3_rsci_radr_d(B_3_rsci_radr_d),
      .B_3_rsci_re_d(B_3_rsci_re_d),
      .B_3_rsci_q_d(B_3_rsci_q_d),
      .P_W_rsci_radr_d(P_W_rsci_radr_d),
      .P_W_rsci_re_d(P_W_rsci_re_d),
      .P_W_rsci_q_d(P_W_rsci_q_d),
      .P_B_rsci_radr_d(P_B_rsci_radr_d),
      .P_B_rsci_re_d(P_B_rsci_re_d),
      .P_B_rsci_q_d(P_B_rsci_q_d),
      .memory_1_rsci_radr_d(memory_1_rsci_radr_d),
      .memory_1_rsci_wadr_d(memory_1_rsci_wadr_d),
      .memory_1_rsci_d_d(memory_1_rsci_d_d),
      .memory_1_rsci_we_d(memory_1_rsci_we_d),
      .memory_1_rsci_re_d(memory_1_rsci_re_d),
      .memory_1_rsci_q_d(memory_1_rsci_q_d),
      .memory_2_rsci_radr_d(memory_2_rsci_radr_d),
      .memory_2_rsci_wadr_d(memory_2_rsci_wadr_d),
      .memory_2_rsci_d_d(memory_2_rsci_d_d),
      .memory_2_rsci_we_d(memory_2_rsci_we_d),
      .memory_2_rsci_re_d(memory_2_rsci_re_d),
      .memory_2_rsci_q_d(memory_2_rsci_q_d),
      .image_rsci_re_d_pff(image_rsci_re_d_iff)
    );
endmodule



