
--------> /softl3/catapultc10_1b/Mgc_home/pkgs/siflibs/ccs_out_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_out_pkg_v1 IS

COMPONENT ccs_out_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    dat    : OUT std_logic_vector(width-1 DOWNTO 0);
    idat   : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END ccs_out_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_out_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    dat   : OUT std_logic_vector(width-1 DOWNTO 0);
    idat  : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END ccs_out_v1;

ARCHITECTURE beh OF ccs_out_v1 IS
BEGIN

  dat <= idat;

END beh;


--------> /softl3/catapultc10_1b/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_io_sync_pkg_v2 IS

COMPONENT mgc_io_sync_v2
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END COMPONENT;

END mgc_io_sync_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_io_sync_v2 IS
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END mgc_io_sync_v2;

ARCHITECTURE beh OF mgc_io_sync_v2 IS
BEGIN

  lz <= ld;

END beh;


--------> /softl3/catapultc10_1b/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.vhd 

LIBRARY IEEE;

   USE IEEE.STD_LOGIC_1164.ALL;
   USE IEEE.Numeric_Std.ALL;

PACKAGE BLOCK_1R1W_RBW_pkg IS

   COMPONENT BLOCK_1R1W_RBW
      GENERIC (
         data_width    : integer := 8;
         addr_width : integer := 7;
         depth         : integer := 128
      );
      PORT (
         clk  : IN  std_logic;
         radr : IN  std_logic_vector(addr_width-1 DOWNTO 0);
         wadr : IN  std_logic_vector(addr_width-1 DOWNTO 0);
         we   : IN  std_logic;
         re   : IN  std_logic;
         d    : IN  std_logic_vector(data_width-1 DOWNTO 0);
         q    : OUT std_logic_vector(data_width-1  DOWNTO 0)
      );
   END COMPONENT;

END BLOCK_1R1W_RBW_pkg;


LIBRARY IEEE;

   USE IEEE.STD_LOGIC_1164.ALL;
   USE IEEE.Numeric_Std.ALL;

ENTITY BLOCK_1R1W_RBW IS
      GENERIC (
         data_width    : integer := 8;
         addr_width : integer := 7;
         depth         : integer := 128
      );
      PORT (
         clk  : IN  std_logic;
         radr : IN  std_logic_vector(addr_width-1 DOWNTO 0);
         wadr : IN  std_logic_vector(addr_width-1 DOWNTO 0);
         we   : IN  std_logic;
         re   : IN  std_logic;
         d    : IN  std_logic_vector(data_width-1 DOWNTO 0);
         q    : OUT std_logic_vector(data_width-1  DOWNTO 0)
      );
END BLOCK_1R1W_RBW;

ARCHITECTURE rtl OF BLOCK_1R1W_RBW IS

   TYPE ram_t IS ARRAY (depth-1 DOWNTO 0) OF std_logic_vector(data_width-1 DOWNTO 0);
   SIGNAL mem : ram_t := (OTHERS => (OTHERS => '0'));

   ATTRIBUTE ram_style: STRING;
   ATTRIBUTE ram_style OF mem : SIGNAL IS "BLOCK";
   ATTRIBUTE syn_ramstyle: STRING;
   ATTRIBUTE syn_ramstyle OF mem : SIGNAL IS "block_ram";

BEGIN
   PROCESS (clk)
   BEGIN
      IF (rising_edge(clk)) THEN
         IF (we='1') THEN
           mem(to_integer(unsigned(wadr))) <= d;
         END IF;
         IF (re='1') THEN
            q <= mem(to_integer(unsigned(radr))) ; -- read port
         END IF; 
      END IF;
   END PROCESS;
END rtl;


--------> ./rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.1b/747384 Production Release
--  HLS Date:       Wed Nov  1 10:26:06 PDT 2017
-- 
--  Generated by:   xph3sei710@ocaepc56
--  Generated date: Fri Jan 25 10:40:00 2019
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_11_1728_12_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_11_1728_12_gen IS
  PORT(
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
    re : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    we_d : IN STD_LOGIC;
    re_d : IN STD_LOGIC;
    q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
  );
END CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_11_1728_12_gen;

ARCHITECTURE v18 OF CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_11_1728_12_gen
    IS
  -- Default Constants

BEGIN
  -- Default Constant Signal Assignments

  we <= (we_d);
  d <= (d_d);
  wadr <= (wadr_d);
  re <= (re_d);
  q_d <= q;
  radr <= (radr_d);
END v18;

-- ------------------------------------------------------------------
--  Design Unit:    CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_11_1728_11_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_11_1728_11_gen IS
  PORT(
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
    re : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    we_d : IN STD_LOGIC;
    re_d : IN STD_LOGIC;
    q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
  );
END CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_11_1728_11_gen;

ARCHITECTURE v18 OF CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_11_1728_11_gen
    IS
  -- Default Constants

BEGIN
  -- Default Constant Signal Assignments

  we <= (we_d);
  d <= (d_d);
  wadr <= (wadr_d);
  re <= (re_d);
  q_d <= q;
  radr <= (radr_d);
END v18;

-- ------------------------------------------------------------------
--  Design Unit:    CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_4_10_9_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_4_10_9_gen IS
  PORT(
    re : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    re_d : IN STD_LOGIC;
    q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
  );
END CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_4_10_9_gen;

ARCHITECTURE v18 OF CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_4_10_9_gen
    IS
  -- Default Constants

BEGIN
  -- Default Constant Signal Assignments

  re <= (re_d);
  q_d <= q;
  radr <= (radr_d);
END v18;

-- ------------------------------------------------------------------
--  Design Unit:    CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1800_8_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1800_8_gen IS
  PORT(
    re : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
    re_d : IN STD_LOGIC;
    q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
  );
END CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1800_8_gen;

ARCHITECTURE v18 OF CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1800_8_gen
    IS
  -- Default Constants

BEGIN
  -- Default Constant Signal Assignments

  re <= (re_d);
  q_d <= q;
  radr <= (radr_d);
END v18;

-- ------------------------------------------------------------------
--  Design Unit:    CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_5_20_7_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_5_20_7_gen IS
  PORT(
    re : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    re_d : IN STD_LOGIC;
    q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
  );
END CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_5_20_7_gen;

ARCHITECTURE v18 OF CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_5_20_7_gen
    IS
  -- Default Constants

BEGIN
  -- Default Constant Signal Assignments

  re <= (re_d);
  q_d <= q;
  radr <= (radr_d);
END v18;

-- ------------------------------------------------------------------
--  Design Unit:    CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_13_5760_6_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_13_5760_6_gen IS
  PORT(
    re : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
    re_d : IN STD_LOGIC;
    q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
  );
END CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_13_5760_6_gen;

ARCHITECTURE v18 OF CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_13_5760_6_gen
    IS
  -- Default Constants

BEGIN
  -- Default Constant Signal Assignments

  re <= (re_d);
  q_d <= q;
  radr <= (radr_d);
END v18;

-- ------------------------------------------------------------------
--  Design Unit:    CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_5_32_5_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_5_32_5_gen IS
  PORT(
    re : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    re_d : IN STD_LOGIC;
    q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
  );
END CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_5_32_5_gen;

ARCHITECTURE v18 OF CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_5_32_5_gen
    IS
  -- Default Constants

BEGIN
  -- Default Constant Signal Assignments

  re <= (re_d);
  q_d <= q;
  radr <= (radr_d);
END v18;

-- ------------------------------------------------------------------
--  Design Unit:    CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_15_18432_4_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_15_18432_4_gen IS
  PORT(
    re : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (14 DOWNTO 0);
    re_d : IN STD_LOGIC;
    q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
  );
END CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_15_18432_4_gen;

ARCHITECTURE v18 OF CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_15_18432_4_gen
    IS
  -- Default Constants

BEGIN
  -- Default Constant Signal Assignments

  re <= (re_d);
  q_d <= q;
  radr <= (radr_d);
END v18;

-- ------------------------------------------------------------------
--  Design Unit:    CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_6_64_3_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_6_64_3_gen IS
  PORT(
    re : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    re_d : IN STD_LOGIC;
    q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
  );
END CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_6_64_3_gen;

ARCHITECTURE v18 OF CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_6_64_3_gen
    IS
  -- Default Constants

BEGIN
  -- Default Constant Signal Assignments

  re <= (re_d);
  q_d <= q;
  radr <= (radr_d);
END v18;

-- ------------------------------------------------------------------
--  Design Unit:    CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1728_2_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1728_2_gen IS
  PORT(
    re : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
    re_d : IN STD_LOGIC;
    q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
  );
END CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1728_2_gen;

ARCHITECTURE v18 OF CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1728_2_gen
    IS
  -- Default Constants

BEGIN
  -- Default Constant Signal Assignments

  re <= (re_d);
  q_d <= q;
  radr <= (radr_d);
END v18;

-- ------------------------------------------------------------------
--  Design Unit:    CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1728_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1728_1_gen IS
  PORT(
    re : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
    re_d : IN STD_LOGIC;
    q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
  );
END CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1728_1_gen;

ARCHITECTURE v18 OF CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1728_1_gen
    IS
  -- Default Constants

BEGIN
  -- Default Constant Signal Assignments

  re <= (re_d);
  q_d <= q;
  radr <= (radr_d);
END v18;

-- ------------------------------------------------------------------
--  Design Unit:    CNN_main_simple_core_core_fsm
--  FSM Module
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY CNN_main_simple_core_core_fsm IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    fsm_output : OUT STD_LOGIC_VECTOR (91 DOWNTO 0);
    INIT_I_C_1_tr0 : IN STD_LOGIC;
    INIT_J_C_0_tr0 : IN STD_LOGIC;
    INIT_L_C_0_tr0 : IN STD_LOGIC;
    FOR_B_C_1_tr0 : IN STD_LOGIC;
    FOR_A_C_0_tr0 : IN STD_LOGIC;
    FOR_I_C_2_tr0 : IN STD_LOGIC;
    FOR_J_C_0_tr0 : IN STD_LOGIC;
    FOR_K_C_0_tr0 : IN STD_LOGIC;
    BIAS_I_C_2_tr0 : IN STD_LOGIC;
    BIAS_J_C_0_tr0 : IN STD_LOGIC;
    FOR_L_C_0_tr0 : IN STD_LOGIC;
    FOR_A_1_C_1_tr0 : IN STD_LOGIC;
    FOR_B_1_C_1_tr0 : IN STD_LOGIC;
    FOR_I_1_C_1_tr0 : IN STD_LOGIC;
    FOR_J_1_C_1_tr0 : IN STD_LOGIC;
    FOR_K_1_C_0_tr0 : IN STD_LOGIC;
    INIT_I_1_C_1_tr0 : IN STD_LOGIC;
    INIT_J_1_C_0_tr0 : IN STD_LOGIC;
    INIT_L_1_C_0_tr0 : IN STD_LOGIC;
    FOR_B_2_C_1_tr0 : IN STD_LOGIC;
    FOR_A_2_C_0_tr0 : IN STD_LOGIC;
    FOR_I_2_C_2_tr0 : IN STD_LOGIC;
    FOR_J_2_C_0_tr0 : IN STD_LOGIC;
    FOR_K_2_C_0_tr0 : IN STD_LOGIC;
    BIAS_I_1_C_2_tr0 : IN STD_LOGIC;
    BIAS_J_1_C_0_tr0 : IN STD_LOGIC;
    FOR_L_1_C_0_tr0 : IN STD_LOGIC;
    FOR_A_3_C_1_tr0 : IN STD_LOGIC;
    FOR_B_3_C_1_tr0 : IN STD_LOGIC;
    FOR_I_3_C_1_tr0 : IN STD_LOGIC;
    FOR_J_3_C_1_tr0 : IN STD_LOGIC;
    FOR_K_3_C_0_tr0 : IN STD_LOGIC;
    INIT_I_2_C_1_tr0 : IN STD_LOGIC;
    INIT_J_2_C_0_tr0 : IN STD_LOGIC;
    INIT_L_2_C_0_tr0 : IN STD_LOGIC;
    FOR_B_4_C_1_tr0 : IN STD_LOGIC;
    FOR_A_4_C_0_tr0 : IN STD_LOGIC;
    FOR_I_4_C_2_tr0 : IN STD_LOGIC;
    FOR_J_4_C_0_tr0 : IN STD_LOGIC;
    FOR_K_4_C_0_tr0 : IN STD_LOGIC;
    BIAS_I_2_C_2_tr0 : IN STD_LOGIC;
    BIAS_J_2_C_0_tr0 : IN STD_LOGIC;
    FOR_L_2_C_0_tr0 : IN STD_LOGIC;
    FOR_A_5_C_1_tr0 : IN STD_LOGIC;
    FOR_B_5_C_1_tr0 : IN STD_LOGIC;
    FOR_I_5_C_1_tr0 : IN STD_LOGIC;
    FOR_J_5_C_1_tr0 : IN STD_LOGIC;
    FOR_K_5_C_0_tr0 : IN STD_LOGIC;
    FOR_K_6_C_2_tr0 : IN STD_LOGIC;
    FOR_J_6_C_0_tr0 : IN STD_LOGIC;
    FOR_I_6_C_0_tr0 : IN STD_LOGIC;
    FOR_K_7_C_1_tr0 : IN STD_LOGIC;
    FOR_J_7_C_1_tr0 : IN STD_LOGIC;
    for_C_0_tr0 : IN STD_LOGIC
  );
END CNN_main_simple_core_core_fsm;

ARCHITECTURE v18 OF CNN_main_simple_core_core_fsm IS
  -- Default Constants

  -- FSM State Type Declaration for CNN_main_simple_core_core_fsm_1
  TYPE CNN_main_simple_core_core_fsm_1_ST IS (core_rlp_C_0, core_rlp_C_1, main_C_0,
      INIT_I_C_0, INIT_I_C_1, INIT_J_C_0, INIT_L_C_0, FOR_B_C_0, FOR_B_C_1, FOR_A_C_0,
      FOR_I_C_0, FOR_I_C_1, FOR_I_C_2, FOR_J_C_0, FOR_K_C_0, BIAS_I_C_0, BIAS_I_C_1,
      BIAS_I_C_2, BIAS_J_C_0, FOR_L_C_0, FOR_J_1_C_0, FOR_I_1_C_0, FOR_A_1_C_0, FOR_A_1_C_1,
      FOR_B_1_C_0, FOR_B_1_C_1, FOR_I_1_C_1, FOR_J_1_C_1, FOR_K_1_C_0, INIT_I_1_C_0,
      INIT_I_1_C_1, INIT_J_1_C_0, INIT_L_1_C_0, FOR_B_2_C_0, FOR_B_2_C_1, FOR_A_2_C_0,
      FOR_I_2_C_0, FOR_I_2_C_1, FOR_I_2_C_2, FOR_J_2_C_0, FOR_K_2_C_0, BIAS_I_1_C_0,
      BIAS_I_1_C_1, BIAS_I_1_C_2, BIAS_J_1_C_0, FOR_L_1_C_0, FOR_J_3_C_0, FOR_I_3_C_0,
      FOR_A_3_C_0, FOR_A_3_C_1, FOR_B_3_C_0, FOR_B_3_C_1, FOR_I_3_C_1, FOR_J_3_C_1,
      FOR_K_3_C_0, INIT_I_2_C_0, INIT_I_2_C_1, INIT_J_2_C_0, INIT_L_2_C_0, FOR_B_4_C_0,
      FOR_B_4_C_1, FOR_A_4_C_0, FOR_I_4_C_0, FOR_I_4_C_1, FOR_I_4_C_2, FOR_J_4_C_0,
      FOR_K_4_C_0, BIAS_I_2_C_0, BIAS_I_2_C_1, BIAS_I_2_C_2, BIAS_J_2_C_0, FOR_L_2_C_0,
      FOR_J_5_C_0, FOR_I_5_C_0, FOR_A_5_C_0, FOR_A_5_C_1, FOR_B_5_C_0, FOR_B_5_C_1,
      FOR_I_5_C_1, FOR_J_5_C_1, FOR_K_5_C_0, FOR_K_6_C_0, FOR_K_6_C_1, FOR_K_6_C_2,
      FOR_J_6_C_0, FOR_I_6_C_0, FOR_J_7_C_0, FOR_K_7_C_0, FOR_K_7_C_1, FOR_J_7_C_1,
      for_C_0, main_C_1);

  SIGNAL state_var : CNN_main_simple_core_core_fsm_1_ST;
  SIGNAL state_var_NS : CNN_main_simple_core_core_fsm_1_ST;

BEGIN
  -- Default Constant Signal Assignments

  CNN_main_simple_core_core_fsm_1 : PROCESS (INIT_I_C_1_tr0, INIT_J_C_0_tr0, INIT_L_C_0_tr0,
      FOR_B_C_1_tr0, FOR_A_C_0_tr0, FOR_I_C_2_tr0, FOR_J_C_0_tr0, FOR_K_C_0_tr0,
      BIAS_I_C_2_tr0, BIAS_J_C_0_tr0, FOR_L_C_0_tr0, FOR_A_1_C_1_tr0, FOR_B_1_C_1_tr0,
      FOR_I_1_C_1_tr0, FOR_J_1_C_1_tr0, FOR_K_1_C_0_tr0, INIT_I_1_C_1_tr0, INIT_J_1_C_0_tr0,
      INIT_L_1_C_0_tr0, FOR_B_2_C_1_tr0, FOR_A_2_C_0_tr0, FOR_I_2_C_2_tr0, FOR_J_2_C_0_tr0,
      FOR_K_2_C_0_tr0, BIAS_I_1_C_2_tr0, BIAS_J_1_C_0_tr0, FOR_L_1_C_0_tr0, FOR_A_3_C_1_tr0,
      FOR_B_3_C_1_tr0, FOR_I_3_C_1_tr0, FOR_J_3_C_1_tr0, FOR_K_3_C_0_tr0, INIT_I_2_C_1_tr0,
      INIT_J_2_C_0_tr0, INIT_L_2_C_0_tr0, FOR_B_4_C_1_tr0, FOR_A_4_C_0_tr0, FOR_I_4_C_2_tr0,
      FOR_J_4_C_0_tr0, FOR_K_4_C_0_tr0, BIAS_I_2_C_2_tr0, BIAS_J_2_C_0_tr0, FOR_L_2_C_0_tr0,
      FOR_A_5_C_1_tr0, FOR_B_5_C_1_tr0, FOR_I_5_C_1_tr0, FOR_J_5_C_1_tr0, FOR_K_5_C_0_tr0,
      FOR_K_6_C_2_tr0, FOR_J_6_C_0_tr0, FOR_I_6_C_0_tr0, FOR_K_7_C_1_tr0, FOR_J_7_C_1_tr0,
      for_C_0_tr0, state_var)
  BEGIN
    CASE state_var IS
      WHEN core_rlp_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010");
        state_var_NS <= main_C_0;
      WHEN main_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100");
        state_var_NS <= INIT_I_C_0;
      WHEN INIT_I_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000");
        state_var_NS <= INIT_I_C_1;
      WHEN INIT_I_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000");
        IF ( INIT_I_C_1_tr0 = '1' ) THEN
          state_var_NS <= INIT_J_C_0;
        ELSE
          state_var_NS <= INIT_I_C_0;
        END IF;
      WHEN INIT_J_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000");
        IF ( INIT_J_C_0_tr0 = '1' ) THEN
          state_var_NS <= INIT_L_C_0;
        ELSE
          state_var_NS <= INIT_I_C_0;
        END IF;
      WHEN INIT_L_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000");
        IF ( INIT_L_C_0_tr0 = '1' ) THEN
          state_var_NS <= FOR_B_C_0;
        ELSE
          state_var_NS <= INIT_I_C_0;
        END IF;
      WHEN FOR_B_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000");
        state_var_NS <= FOR_B_C_1;
      WHEN FOR_B_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000");
        IF ( FOR_B_C_1_tr0 = '1' ) THEN
          state_var_NS <= FOR_A_C_0;
        ELSE
          state_var_NS <= FOR_B_C_0;
        END IF;
      WHEN FOR_A_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000");
        IF ( FOR_A_C_0_tr0 = '1' ) THEN
          state_var_NS <= FOR_I_C_0;
        ELSE
          state_var_NS <= FOR_B_C_0;
        END IF;
      WHEN FOR_I_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000");
        state_var_NS <= FOR_I_C_1;
      WHEN FOR_I_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000");
        state_var_NS <= FOR_I_C_2;
      WHEN FOR_I_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000");
        IF ( FOR_I_C_2_tr0 = '1' ) THEN
          state_var_NS <= FOR_J_C_0;
        ELSE
          state_var_NS <= FOR_B_C_0;
        END IF;
      WHEN FOR_J_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000");
        IF ( FOR_J_C_0_tr0 = '1' ) THEN
          state_var_NS <= FOR_K_C_0;
        ELSE
          state_var_NS <= FOR_B_C_0;
        END IF;
      WHEN FOR_K_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000");
        IF ( FOR_K_C_0_tr0 = '1' ) THEN
          state_var_NS <= BIAS_I_C_0;
        ELSE
          state_var_NS <= FOR_B_C_0;
        END IF;
      WHEN BIAS_I_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000");
        state_var_NS <= BIAS_I_C_1;
      WHEN BIAS_I_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000");
        state_var_NS <= BIAS_I_C_2;
      WHEN BIAS_I_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000");
        IF ( BIAS_I_C_2_tr0 = '1' ) THEN
          state_var_NS <= BIAS_J_C_0;
        ELSE
          state_var_NS <= BIAS_I_C_0;
        END IF;
      WHEN BIAS_J_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000");
        IF ( BIAS_J_C_0_tr0 = '1' ) THEN
          state_var_NS <= FOR_L_C_0;
        ELSE
          state_var_NS <= BIAS_I_C_0;
        END IF;
      WHEN FOR_L_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000");
        IF ( FOR_L_C_0_tr0 = '1' ) THEN
          state_var_NS <= FOR_J_1_C_0;
        ELSE
          state_var_NS <= FOR_B_C_0;
        END IF;
      WHEN FOR_J_1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000");
        state_var_NS <= FOR_I_1_C_0;
      WHEN FOR_I_1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000");
        state_var_NS <= FOR_A_1_C_0;
      WHEN FOR_A_1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000");
        state_var_NS <= FOR_A_1_C_1;
      WHEN FOR_A_1_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000");
        IF ( FOR_A_1_C_1_tr0 = '1' ) THEN
          state_var_NS <= FOR_B_1_C_0;
        ELSE
          state_var_NS <= FOR_A_1_C_0;
        END IF;
      WHEN FOR_B_1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000");
        state_var_NS <= FOR_B_1_C_1;
      WHEN FOR_B_1_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000");
        IF ( FOR_B_1_C_1_tr0 = '1' ) THEN
          state_var_NS <= FOR_I_1_C_1;
        ELSE
          state_var_NS <= FOR_A_1_C_0;
        END IF;
      WHEN FOR_I_1_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000");
        IF ( FOR_I_1_C_1_tr0 = '1' ) THEN
          state_var_NS <= FOR_J_1_C_1;
        ELSE
          state_var_NS <= FOR_I_1_C_0;
        END IF;
      WHEN FOR_J_1_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000");
        IF ( FOR_J_1_C_1_tr0 = '1' ) THEN
          state_var_NS <= FOR_K_1_C_0;
        ELSE
          state_var_NS <= FOR_J_1_C_0;
        END IF;
      WHEN FOR_K_1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000");
        IF ( FOR_K_1_C_0_tr0 = '1' ) THEN
          state_var_NS <= INIT_I_1_C_0;
        ELSE
          state_var_NS <= FOR_J_1_C_0;
        END IF;
      WHEN INIT_I_1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000");
        state_var_NS <= INIT_I_1_C_1;
      WHEN INIT_I_1_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000");
        IF ( INIT_I_1_C_1_tr0 = '1' ) THEN
          state_var_NS <= INIT_J_1_C_0;
        ELSE
          state_var_NS <= INIT_I_1_C_0;
        END IF;
      WHEN INIT_J_1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000");
        IF ( INIT_J_1_C_0_tr0 = '1' ) THEN
          state_var_NS <= INIT_L_1_C_0;
        ELSE
          state_var_NS <= INIT_I_1_C_0;
        END IF;
      WHEN INIT_L_1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000");
        IF ( INIT_L_1_C_0_tr0 = '1' ) THEN
          state_var_NS <= FOR_B_2_C_0;
        ELSE
          state_var_NS <= INIT_I_1_C_0;
        END IF;
      WHEN FOR_B_2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000");
        state_var_NS <= FOR_B_2_C_1;
      WHEN FOR_B_2_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000");
        IF ( FOR_B_2_C_1_tr0 = '1' ) THEN
          state_var_NS <= FOR_A_2_C_0;
        ELSE
          state_var_NS <= FOR_B_2_C_0;
        END IF;
      WHEN FOR_A_2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000");
        IF ( FOR_A_2_C_0_tr0 = '1' ) THEN
          state_var_NS <= FOR_I_2_C_0;
        ELSE
          state_var_NS <= FOR_B_2_C_0;
        END IF;
      WHEN FOR_I_2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000");
        state_var_NS <= FOR_I_2_C_1;
      WHEN FOR_I_2_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000");
        state_var_NS <= FOR_I_2_C_2;
      WHEN FOR_I_2_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000");
        IF ( FOR_I_2_C_2_tr0 = '1' ) THEN
          state_var_NS <= FOR_J_2_C_0;
        ELSE
          state_var_NS <= FOR_B_2_C_0;
        END IF;
      WHEN FOR_J_2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000");
        IF ( FOR_J_2_C_0_tr0 = '1' ) THEN
          state_var_NS <= FOR_K_2_C_0;
        ELSE
          state_var_NS <= FOR_B_2_C_0;
        END IF;
      WHEN FOR_K_2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000");
        IF ( FOR_K_2_C_0_tr0 = '1' ) THEN
          state_var_NS <= BIAS_I_1_C_0;
        ELSE
          state_var_NS <= FOR_B_2_C_0;
        END IF;
      WHEN BIAS_I_1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000");
        state_var_NS <= BIAS_I_1_C_1;
      WHEN BIAS_I_1_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000");
        state_var_NS <= BIAS_I_1_C_2;
      WHEN BIAS_I_1_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000");
        IF ( BIAS_I_1_C_2_tr0 = '1' ) THEN
          state_var_NS <= BIAS_J_1_C_0;
        ELSE
          state_var_NS <= BIAS_I_1_C_0;
        END IF;
      WHEN BIAS_J_1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000");
        IF ( BIAS_J_1_C_0_tr0 = '1' ) THEN
          state_var_NS <= FOR_L_1_C_0;
        ELSE
          state_var_NS <= BIAS_I_1_C_0;
        END IF;
      WHEN FOR_L_1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000");
        IF ( FOR_L_1_C_0_tr0 = '1' ) THEN
          state_var_NS <= FOR_J_3_C_0;
        ELSE
          state_var_NS <= FOR_B_2_C_0;
        END IF;
      WHEN FOR_J_3_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000");
        state_var_NS <= FOR_I_3_C_0;
      WHEN FOR_I_3_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000");
        state_var_NS <= FOR_A_3_C_0;
      WHEN FOR_A_3_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000");
        state_var_NS <= FOR_A_3_C_1;
      WHEN FOR_A_3_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000");
        IF ( FOR_A_3_C_1_tr0 = '1' ) THEN
          state_var_NS <= FOR_B_3_C_0;
        ELSE
          state_var_NS <= FOR_A_3_C_0;
        END IF;
      WHEN FOR_B_3_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000");
        state_var_NS <= FOR_B_3_C_1;
      WHEN FOR_B_3_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000");
        IF ( FOR_B_3_C_1_tr0 = '1' ) THEN
          state_var_NS <= FOR_I_3_C_1;
        ELSE
          state_var_NS <= FOR_A_3_C_0;
        END IF;
      WHEN FOR_I_3_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000");
        IF ( FOR_I_3_C_1_tr0 = '1' ) THEN
          state_var_NS <= FOR_J_3_C_1;
        ELSE
          state_var_NS <= FOR_I_3_C_0;
        END IF;
      WHEN FOR_J_3_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000");
        IF ( FOR_J_3_C_1_tr0 = '1' ) THEN
          state_var_NS <= FOR_K_3_C_0;
        ELSE
          state_var_NS <= FOR_J_3_C_0;
        END IF;
      WHEN FOR_K_3_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000");
        IF ( FOR_K_3_C_0_tr0 = '1' ) THEN
          state_var_NS <= INIT_I_2_C_0;
        ELSE
          state_var_NS <= FOR_J_3_C_0;
        END IF;
      WHEN INIT_I_2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000");
        state_var_NS <= INIT_I_2_C_1;
      WHEN INIT_I_2_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000");
        IF ( INIT_I_2_C_1_tr0 = '1' ) THEN
          state_var_NS <= INIT_J_2_C_0;
        ELSE
          state_var_NS <= INIT_I_2_C_0;
        END IF;
      WHEN INIT_J_2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000");
        IF ( INIT_J_2_C_0_tr0 = '1' ) THEN
          state_var_NS <= INIT_L_2_C_0;
        ELSE
          state_var_NS <= INIT_I_2_C_0;
        END IF;
      WHEN INIT_L_2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000");
        IF ( INIT_L_2_C_0_tr0 = '1' ) THEN
          state_var_NS <= FOR_B_4_C_0;
        ELSE
          state_var_NS <= INIT_I_2_C_0;
        END IF;
      WHEN FOR_B_4_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000");
        state_var_NS <= FOR_B_4_C_1;
      WHEN FOR_B_4_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000");
        IF ( FOR_B_4_C_1_tr0 = '1' ) THEN
          state_var_NS <= FOR_A_4_C_0;
        ELSE
          state_var_NS <= FOR_B_4_C_0;
        END IF;
      WHEN FOR_A_4_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000");
        IF ( FOR_A_4_C_0_tr0 = '1' ) THEN
          state_var_NS <= FOR_I_4_C_0;
        ELSE
          state_var_NS <= FOR_B_4_C_0;
        END IF;
      WHEN FOR_I_4_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000");
        state_var_NS <= FOR_I_4_C_1;
      WHEN FOR_I_4_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000");
        state_var_NS <= FOR_I_4_C_2;
      WHEN FOR_I_4_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000");
        IF ( FOR_I_4_C_2_tr0 = '1' ) THEN
          state_var_NS <= FOR_J_4_C_0;
        ELSE
          state_var_NS <= FOR_B_4_C_0;
        END IF;
      WHEN FOR_J_4_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000");
        IF ( FOR_J_4_C_0_tr0 = '1' ) THEN
          state_var_NS <= FOR_K_4_C_0;
        ELSE
          state_var_NS <= FOR_B_4_C_0;
        END IF;
      WHEN FOR_K_4_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000");
        IF ( FOR_K_4_C_0_tr0 = '1' ) THEN
          state_var_NS <= BIAS_I_2_C_0;
        ELSE
          state_var_NS <= FOR_B_4_C_0;
        END IF;
      WHEN BIAS_I_2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000");
        state_var_NS <= BIAS_I_2_C_1;
      WHEN BIAS_I_2_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000");
        state_var_NS <= BIAS_I_2_C_2;
      WHEN BIAS_I_2_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000");
        IF ( BIAS_I_2_C_2_tr0 = '1' ) THEN
          state_var_NS <= BIAS_J_2_C_0;
        ELSE
          state_var_NS <= BIAS_I_2_C_0;
        END IF;
      WHEN BIAS_J_2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000");
        IF ( BIAS_J_2_C_0_tr0 = '1' ) THEN
          state_var_NS <= FOR_L_2_C_0;
        ELSE
          state_var_NS <= BIAS_I_2_C_0;
        END IF;
      WHEN FOR_L_2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000");
        IF ( FOR_L_2_C_0_tr0 = '1' ) THEN
          state_var_NS <= FOR_J_5_C_0;
        ELSE
          state_var_NS <= FOR_B_4_C_0;
        END IF;
      WHEN FOR_J_5_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000");
        state_var_NS <= FOR_I_5_C_0;
      WHEN FOR_I_5_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000");
        state_var_NS <= FOR_A_5_C_0;
      WHEN FOR_A_5_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000");
        state_var_NS <= FOR_A_5_C_1;
      WHEN FOR_A_5_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000");
        IF ( FOR_A_5_C_1_tr0 = '1' ) THEN
          state_var_NS <= FOR_B_5_C_0;
        ELSE
          state_var_NS <= FOR_A_5_C_0;
        END IF;
      WHEN FOR_B_5_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000");
        state_var_NS <= FOR_B_5_C_1;
      WHEN FOR_B_5_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000");
        IF ( FOR_B_5_C_1_tr0 = '1' ) THEN
          state_var_NS <= FOR_I_5_C_1;
        ELSE
          state_var_NS <= FOR_A_5_C_0;
        END IF;
      WHEN FOR_I_5_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000");
        IF ( FOR_I_5_C_1_tr0 = '1' ) THEN
          state_var_NS <= FOR_J_5_C_1;
        ELSE
          state_var_NS <= FOR_I_5_C_0;
        END IF;
      WHEN FOR_J_5_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000");
        IF ( FOR_J_5_C_1_tr0 = '1' ) THEN
          state_var_NS <= FOR_K_5_C_0;
        ELSE
          state_var_NS <= FOR_J_5_C_0;
        END IF;
      WHEN FOR_K_5_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000");
        IF ( FOR_K_5_C_0_tr0 = '1' ) THEN
          state_var_NS <= FOR_K_6_C_0;
        ELSE
          state_var_NS <= FOR_J_5_C_0;
        END IF;
      WHEN FOR_K_6_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000");
        state_var_NS <= FOR_K_6_C_1;
      WHEN FOR_K_6_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000");
        state_var_NS <= FOR_K_6_C_2;
      WHEN FOR_K_6_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000");
        IF ( FOR_K_6_C_2_tr0 = '1' ) THEN
          state_var_NS <= FOR_J_6_C_0;
        ELSE
          state_var_NS <= FOR_K_6_C_0;
        END IF;
      WHEN FOR_J_6_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
        IF ( FOR_J_6_C_0_tr0 = '1' ) THEN
          state_var_NS <= FOR_I_6_C_0;
        ELSE
          state_var_NS <= FOR_K_6_C_0;
        END IF;
      WHEN FOR_I_6_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
        IF ( FOR_I_6_C_0_tr0 = '1' ) THEN
          state_var_NS <= FOR_J_7_C_0;
        ELSE
          state_var_NS <= FOR_K_6_C_0;
        END IF;
      WHEN FOR_J_7_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
        state_var_NS <= FOR_K_7_C_0;
      WHEN FOR_K_7_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
        state_var_NS <= FOR_K_7_C_1;
      WHEN FOR_K_7_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
        IF ( FOR_K_7_C_1_tr0 = '1' ) THEN
          state_var_NS <= FOR_J_7_C_1;
        ELSE
          state_var_NS <= FOR_K_7_C_0;
        END IF;
      WHEN FOR_J_7_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
        IF ( FOR_J_7_C_1_tr0 = '1' ) THEN
          state_var_NS <= for_C_0;
        ELSE
          state_var_NS <= FOR_J_7_C_0;
        END IF;
      WHEN for_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
        IF ( for_C_0_tr0 = '1' ) THEN
          state_var_NS <= main_C_1;
        ELSE
          state_var_NS <= for_C_0;
        END IF;
      WHEN main_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
        state_var_NS <= main_C_0;
      -- core_rlp_C_0
      WHEN OTHERS =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001");
        state_var_NS <= core_rlp_C_1;
    END CASE;
  END PROCESS CNN_main_simple_core_core_fsm_1;

  CNN_main_simple_core_core_fsm_1_REG : PROCESS (clk)
  BEGIN
    IF clk'event AND ( clk = '1' ) THEN
      IF ( rst = '1' ) THEN
        state_var <= core_rlp_C_0;
      ELSE
        state_var <= state_var_NS;
      END IF;
    END IF;
  END PROCESS CNN_main_simple_core_core_fsm_1_REG;

END v18;

-- ------------------------------------------------------------------
--  Design Unit:    CNN_main_simple_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY CNN_main_simple_core IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    image_rsc_triosy_lz : OUT STD_LOGIC;
    F_1_rsc_triosy_lz : OUT STD_LOGIC;
    B_1_rsc_triosy_lz : OUT STD_LOGIC;
    F_2_rsc_triosy_lz : OUT STD_LOGIC;
    B_2_rsc_triosy_lz : OUT STD_LOGIC;
    F_3_rsc_triosy_lz : OUT STD_LOGIC;
    B_3_rsc_triosy_lz : OUT STD_LOGIC;
    P_W_rsc_triosy_lz : OUT STD_LOGIC;
    P_B_rsc_triosy_lz : OUT STD_LOGIC;
    index_rsc_dat : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    index_rsc_triosy_lz : OUT STD_LOGIC;
    image_rsci_radr_d : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
    image_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    F_1_rsci_radr_d : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
    F_1_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    B_1_rsci_radr_d : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    B_1_rsci_re_d : OUT STD_LOGIC;
    B_1_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    F_2_rsci_radr_d : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
    F_2_rsci_re_d : OUT STD_LOGIC;
    F_2_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    B_2_rsci_radr_d : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    B_2_rsci_re_d : OUT STD_LOGIC;
    B_2_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    F_3_rsci_radr_d : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
    F_3_rsci_re_d : OUT STD_LOGIC;
    F_3_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    B_3_rsci_radr_d : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    B_3_rsci_re_d : OUT STD_LOGIC;
    B_3_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    P_W_rsci_radr_d : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
    P_W_rsci_re_d : OUT STD_LOGIC;
    P_W_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    P_B_rsci_radr_d : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    P_B_rsci_re_d : OUT STD_LOGIC;
    P_B_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    memory_1_rsci_radr_d : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
    memory_1_rsci_wadr_d : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
    memory_1_rsci_d_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    memory_1_rsci_we_d : OUT STD_LOGIC;
    memory_1_rsci_re_d : OUT STD_LOGIC;
    memory_1_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    memory_2_rsci_radr_d : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
    memory_2_rsci_wadr_d : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
    memory_2_rsci_d_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    memory_2_rsci_we_d : OUT STD_LOGIC;
    memory_2_rsci_re_d : OUT STD_LOGIC;
    memory_2_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    image_rsci_re_d_pff : OUT STD_LOGIC
  );
END CNN_main_simple_core;

ARCHITECTURE v18 OF CNN_main_simple_core IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL index_rsci_idat : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL fsm_output : STD_LOGIC_VECTOR (91 DOWNTO 0);
  SIGNAL or_dcpl_53 : STD_LOGIC;
  SIGNAL and_dcpl_6 : STD_LOGIC;
  SIGNAL and_dcpl_133 : STD_LOGIC;
  SIGNAL or_dcpl_130 : STD_LOGIC;
  SIGNAL or_dcpl_131 : STD_LOGIC;
  SIGNAL and_dcpl_136 : STD_LOGIC;
  SIGNAL or_dcpl_134 : STD_LOGIC;
  SIGNAL or_dcpl_135 : STD_LOGIC;
  SIGNAL and_dcpl_141 : STD_LOGIC;
  SIGNAL or_dcpl_139 : STD_LOGIC;
  SIGNAL or_dcpl_140 : STD_LOGIC;
  SIGNAL or_dcpl_142 : STD_LOGIC;
  SIGNAL or_tmp_111 : STD_LOGIC;
  SIGNAL or_tmp_117 : STD_LOGIC;
  SIGNAL or_tmp_125 : STD_LOGIC;
  SIGNAL or_tmp_376 : STD_LOGIC;
  SIGNAL or_tmp_379 : STD_LOGIC;
  SIGNAL or_tmp_380 : STD_LOGIC;
  SIGNAL or_tmp_383 : STD_LOGIC;
  SIGNAL or_tmp_392 : STD_LOGIC;
  SIGNAL or_tmp_393 : STD_LOGIC;
  SIGNAL or_tmp_405 : STD_LOGIC;
  SIGNAL or_tmp_406 : STD_LOGIC;
  SIGNAL or_tmp_418 : STD_LOGIC;
  SIGNAL or_tmp_419 : STD_LOGIC;
  SIGNAL or_tmp_431 : STD_LOGIC;
  SIGNAL or_tmp_432 : STD_LOGIC;
  SIGNAL or_tmp_444 : STD_LOGIC;
  SIGNAL or_tmp_445 : STD_LOGIC;
  SIGNAL or_tmp_457 : STD_LOGIC;
  SIGNAL or_tmp_458 : STD_LOGIC;
  SIGNAL or_tmp_470 : STD_LOGIC;
  SIGNAL or_tmp_471 : STD_LOGIC;
  SIGNAL or_tmp_483 : STD_LOGIC;
  SIGNAL or_tmp_484 : STD_LOGIC;
  SIGNAL or_tmp_496 : STD_LOGIC;
  SIGNAL or_tmp_497 : STD_LOGIC;
  SIGNAL FOR_B_4_oelse_acc_tmp_15 : STD_LOGIC;
  SIGNAL FOR_B_2_oelse_acc_tmp_14 : STD_LOGIC;
  SIGNAL FOR_B_oelse_acc_tmp_13 : STD_LOGIC;
  SIGNAL and_4_cse : STD_LOGIC;
  SIGNAL and_10_cse : STD_LOGIC;
  SIGNAL and_16_cse : STD_LOGIC;
  SIGNAL and_285_cse : STD_LOGIC;
  SIGNAL and_283_cse : STD_LOGIC;
  SIGNAL and_316_cse : STD_LOGIC;
  SIGNAL and_318_cse : STD_LOGIC;
  SIGNAL and_317_cse : STD_LOGIC;
  SIGNAL and_386_cse : STD_LOGIC;
  SIGNAL and_307_cse : STD_LOGIC;
  SIGNAL FOR_K_7_slc_FOR_K_7_acc_6_itm : STD_LOGIC;
  SIGNAL FOR_K_7_mux_28_itm : STD_LOGIC;
  SIGNAL FOR_K_7_mux_29_itm : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL FOR_K_7_mux_30_itm : STD_LOGIC;
  SIGNAL FOR_J_7_and_stg_2_1_sva_1 : STD_LOGIC;
  SIGNAL FOR_J_7_and_stg_2_0_sva_1 : STD_LOGIC;
  SIGNAL FOR_J_7_and_stg_1_3_sva_1 : STD_LOGIC;
  SIGNAL FOR_J_7_and_stg_1_2_sva_1 : STD_LOGIC;
  SIGNAL FOR_J_7_and_stg_1_1_sva_1 : STD_LOGIC;
  SIGNAL FOR_J_7_and_stg_1_0_sva_1 : STD_LOGIC;
  SIGNAL FOR_K_6_slc_FOR_K_6_acc_3_itm : STD_LOGIC;
  SIGNAL MP3_simple_a_1_0_sva : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL BIAS_I_2_slc_BIAS_I_2_acc_2_itm : STD_LOGIC;
  SIGNAL BIAS_I_2_slc_15_1_itm : STD_LOGIC_VECTOR (14 DOWNTO 0);
  SIGNAL FOR_I_4_slc_FOR_I_4_acc_2_itm : STD_LOGIC;
  SIGNAL CR3_simple_aux_15_lpi_7_dfm : STD_LOGIC;
  SIGNAL CR3_simple_aux_14_1_lpi_7_dfm : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL CR3_simple_aux_0_lpi_7_dfm : STD_LOGIC;
  SIGNAL CR3_simple_aux_15_lpi_7 : STD_LOGIC;
  SIGNAL CR3_simple_aux_14_1_lpi_7 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL CR3_simple_aux_0_lpi_7 : STD_LOGIC;
  SIGNAL BIAS_I_1_slc_BIAS_I_1_acc_2_itm : STD_LOGIC;
  SIGNAL BIAS_I_1_slc_15_1_itm : STD_LOGIC_VECTOR (14 DOWNTO 0);
  SIGNAL FOR_I_2_slc_FOR_I_2_acc_2_itm : STD_LOGIC;
  SIGNAL CR2_simple_aux_15_lpi_7_dfm : STD_LOGIC;
  SIGNAL CR2_simple_aux_14_1_lpi_7_dfm : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL CR2_simple_aux_0_lpi_7_dfm : STD_LOGIC;
  SIGNAL CR2_simple_aux_15_lpi_7 : STD_LOGIC;
  SIGNAL CR2_simple_aux_14_1_lpi_7 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL CR2_simple_aux_0_lpi_7 : STD_LOGIC;
  SIGNAL BIAS_I_slc_BIAS_I_acc_2_itm : STD_LOGIC;
  SIGNAL BIAS_I_slc_15_1_itm : STD_LOGIC_VECTOR (14 DOWNTO 0);
  SIGNAL FOR_I_slc_FOR_I_acc_2_itm : STD_LOGIC;
  SIGNAL CR1_simple_aux_15_lpi_7_dfm : STD_LOGIC;
  SIGNAL CR1_simple_aux_14_1_lpi_7_dfm : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL CR1_simple_aux_0_lpi_7_dfm : STD_LOGIC;
  SIGNAL CR1_simple_aux_15_lpi_7 : STD_LOGIC;
  SIGNAL CR1_simple_aux_14_1_lpi_7 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL CR1_simple_aux_0_lpi_7 : STD_LOGIC;
  SIGNAL FOR_J_7_and_21_cse_sva : STD_LOGIC;
  SIGNAL FOR_J_7_and_20_cse_sva : STD_LOGIC;
  SIGNAL FOR_J_7_and_19_cse_sva : STD_LOGIC;
  SIGNAL FOR_J_7_and_18_cse_sva : STD_LOGIC;
  SIGNAL FOR_J_7_and_17_cse_sva : STD_LOGIC;
  SIGNAL FOR_J_7_and_16_cse_sva : STD_LOGIC;
  SIGNAL FOR_J_7_and_15_cse_sva : STD_LOGIC;
  SIGNAL FOR_J_7_and_14_cse_sva : STD_LOGIC;
  SIGNAL FOR_J_7_and_13_cse_sva : STD_LOGIC;
  SIGNAL FOR_J_7_and_12_cse_sva : STD_LOGIC;
  SIGNAL perceptron_simple_j_3_0_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL max_sva_15 : STD_LOGIC;
  SIGNAL max_sva_14_1 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL max_sva_0 : STD_LOGIC;
  SIGNAL for_slc_Prob_16_15_0_cse_sva_15_1 : STD_LOGIC;
  SIGNAL for_slc_Prob_16_15_0_cse_sva_14_1_1 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL for_slc_Prob_16_15_0_cse_sva_0_1 : STD_LOGIC;
  SIGNAL MP3_simple_bigger_lpi_6 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL MP2_simple_bigger_lpi_6 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL MP1_simple_bigger_lpi_6 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL CR1_simple_b_1_0_sva_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL FOR_K_7_acc_7_psp_sva_1 : STD_LOGIC_VECTOR (16 DOWNTO 0);
  SIGNAL FOR_B_if_acc_psp_sva_1 : STD_LOGIC_VECTOR (18 DOWNTO 0);
  SIGNAL FOR_A_1_if_asn_MP1_simple_add_M_10_FOR_A_1_if_acc_sdt : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL INIT_I_asn_CR1_simple_add_AF_10_INIT_I_acc_sdt : STD_LOGIC_VECTOR (4 DOWNTO
      0);
  SIGNAL or_220_ssc : STD_LOGIC;
  SIGNAL FOR_B_4_if_acc_10_sdt_4_0_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL reg_index_rsc_triosy_obj_ld_cse : STD_LOGIC;
  SIGNAL reg_CR1_simple_CR1_simple_aux_or_1_cse : STD_LOGIC;
  SIGNAL or_125_cse : STD_LOGIC;
  SIGNAL reg_CR2_simple_CR2_simple_aux_or_1_cse : STD_LOGIC;
  SIGNAL reg_CR3_simple_CR3_simple_aux_or_1_cse : STD_LOGIC;
  SIGNAL FOR_B_2_if_FOR_B_2_if_or_cse : STD_LOGIC;
  SIGNAL or_332_cse : STD_LOGIC;
  SIGNAL or_400_cse : STD_LOGIC;
  SIGNAL or_468_cse : STD_LOGIC;
  SIGNAL FOR_B_4_if_FOR_B_4_if_or_cse : STD_LOGIC;
  SIGNAL reg_CR1_simple_l_1_6_0_sva_5_CR1_simple_l_or_cse : STD_LOGIC;
  SIGNAL reg_MP3_simple_b_1_MP3_simple_b_or_cse : STD_LOGIC;
  SIGNAL memory_1_nor_1_seb : STD_LOGIC;
  SIGNAL memory_1_or_1_seb : STD_LOGIC;
  SIGNAL memory_1_or_seb : STD_LOGIC;
  SIGNAL FOR_K_7_acc_8_sdt_1 : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL perceptron_simple_k_7_0_sva : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL CR3_simple_l_4_0_sva : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL CR2_simple_a_1_0_sva : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL CR2_simple_k_6_0_sva_5_0_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL CR2_simple_l_5_0_sva_4_0_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL CR1_simple_l_6_0_sva_5_0_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL CR1_simple_k_1_0_sva : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL FOR_B_if_acc_10_psp_1 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL FOR_B_if_acc_5_sdt_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL FOR_B_2_if_acc_8_sdt_1 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL FOR_B_2_if_acc_9_psp_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL FOR_B_4_if_acc_11_sdt_1 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL CR3_simple_k_5_0_sva_4_0 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL reshape_simple_k_4_0_sva : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL memory_2_rsci_radr_d_mx0c0 : STD_LOGIC;
  SIGNAL CR2_simple_j_aux_4_0_sva_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL FOR_B_4_if_acc_6_sdt_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL CR3_simple_j_aux_3_0_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL FOR_B_1_if_acc_3_sdt_1 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL MP1_simple_k_6_0_sva_5_0 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL MP2_simple_k_5_0_sva_4_0 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL MP3_simple_k_4_0_sva : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL memory_2_rsci_wadr_d_mx0c0 : STD_LOGIC;
  SIGNAL MP1_simple_i_N_3_0_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL FOR_B_3_if_acc_sdt_1 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL MP2_simple_i_N_2_0_sva_1 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL CR3_simple_a_1_0_sva : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL CR1_simple_a_1_0_sva : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL MP1_simple_bigger_lpi_6_dfm_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL MP2_simple_bigger_lpi_6_dfm_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL MP3_simple_bigger_lpi_6_dfm_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL CR1_simple_j_2_4_0_sva : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL CR1_simple_j_4_0_sva : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL FOR_A_1_oelse_acc_1_ncse_sva_2 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL CR2_simple_j_2_3_0_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL CR2_simple_j_3_0_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL FOR_A_3_oelse_acc_1_ncse_sva_2 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL MP1_simple_a_1_0_sva : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL MP2_simple_a_1_0_sva : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL CR3_simple_j_2_2_0_sva : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL CR3_simple_j_2_0_sva : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL reshape_simple_add_N_10_0_lpi_4 : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL INIT_I_2_acc_6_sdt_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL CR3_simple_l_1_4_0_sva : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL CR1_simple_j_1_4_0_sva : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL CR2_simple_j_1_3_0_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL CR3_simple_j_1_2_0_sva : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL z_out : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL z_out_2 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL z_out_3 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL z_out_4 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL z_out_5 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL z_out_6 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL z_out_7 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL z_out_8 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL z_out_9 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL z_out_10 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL z_out_11 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL z_out_12 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL z_out_13 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL z_out_16 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL z_out_17 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL z_out_19 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL z_out_20 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL z_out_21 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL z_out_22 : STD_LOGIC_VECTOR (16 DOWNTO 0);
  SIGNAL z_out_23 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL z_out_24 : STD_LOGIC_VECTOR (19 DOWNTO 0);
  SIGNAL z_out_25 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL z_out_26 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL CR1_simple_i_1_4_0_sva : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL CR1_simple_i_1_4_0_sva_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL CR1_simple_i_2_4_0_sva : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL CR1_simple_b_1_0_sva : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL CR1_simple_i_2_4_0_sva_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL CR1_simple_i_4_0_sva : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL CR1_simple_i_4_0_sva_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL MP1_simple_j_N_3_0_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL MP1_simple_j_4_1_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL MP1_simple_j_N_3_0_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL MP1_simple_i_N_3_0_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL MP1_simple_i_4_1_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL MP1_simple_b_1_0_sva : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL CR2_simple_i_1_3_0_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL CR2_simple_i_1_3_0_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL CR2_simple_i_2_3_0_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL CR2_simple_b_1_0_sva : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL CR2_simple_i_2_3_0_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL CR2_simple_i_3_0_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL CR2_simple_i_3_0_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL MP2_simple_j_N_2_0_sva : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL MP2_simple_j_3_1_sva : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL MP2_simple_j_N_2_0_sva_1 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL MP2_simple_i_N_2_0_sva : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL MP2_simple_i_3_1_sva : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL MP2_simple_b_1_0_sva : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL CR3_simple_i_1_2_0_sva : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL CR3_simple_i_1_2_0_sva_1 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL CR3_simple_i_2_2_0_sva : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL CR3_simple_b_1_0_sva : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL CR3_simple_i_2_2_0_sva_1 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL CR3_simple_i_2_0_sva : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL CR3_simple_i_2_0_sva_1 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL MP3_simple_j_2_1_sva : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL MP3_simple_j_N_1_0_sva_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL MP3_simple_i_2_1_sva : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL MP3_simple_i_N_1_0_sva_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL MP3_simple_b_1_0_sva : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL reshape_simple_i_1_0_sva : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL reshape_simple_j_1_0_sva : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL reshape_simple_add_N_10_0_sva_1 : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL reshape_simple_k_4_0_sva_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL Prob_4_14_1_sva_1 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL Prob_4_0_sva_1 : STD_LOGIC;
  SIGNAL Prob_4_15_sva_1 : STD_LOGIC;
  SIGNAL Prob_5_14_1_sva_1 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL Prob_5_0_sva_1 : STD_LOGIC;
  SIGNAL Prob_5_15_sva_1 : STD_LOGIC;
  SIGNAL Prob_3_14_1_sva_1 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL Prob_3_0_sva_1 : STD_LOGIC;
  SIGNAL Prob_3_15_sva_1 : STD_LOGIC;
  SIGNAL Prob_6_14_1_sva_1 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL Prob_6_0_sva_1 : STD_LOGIC;
  SIGNAL Prob_6_15_sva_1 : STD_LOGIC;
  SIGNAL Prob_2_14_1_sva_1 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL Prob_2_0_sva_1 : STD_LOGIC;
  SIGNAL Prob_2_15_sva_1 : STD_LOGIC;
  SIGNAL Prob_7_14_1_sva_1 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL Prob_7_0_sva_1 : STD_LOGIC;
  SIGNAL Prob_7_15_sva_1 : STD_LOGIC;
  SIGNAL Prob_1_14_1_sva_1 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL Prob_1_0_sva_1 : STD_LOGIC;
  SIGNAL Prob_1_15_sva_1 : STD_LOGIC;
  SIGNAL Prob_8_14_1_sva_1 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL Prob_8_0_sva_1 : STD_LOGIC;
  SIGNAL Prob_8_15_sva_1 : STD_LOGIC;
  SIGNAL Prob_9_14_1_sva_1 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL Prob_9_0_sva_1 : STD_LOGIC;
  SIGNAL Prob_9_15_sva_1 : STD_LOGIC;
  SIGNAL Prob_4_14_1_sva_2 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL Prob_4_0_sva_2 : STD_LOGIC;
  SIGNAL Prob_4_15_sva_2 : STD_LOGIC;
  SIGNAL Prob_5_14_1_sva_2 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL Prob_5_0_sva_2 : STD_LOGIC;
  SIGNAL Prob_5_15_sva_2 : STD_LOGIC;
  SIGNAL Prob_3_14_1_sva_2 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL Prob_3_0_sva_2 : STD_LOGIC;
  SIGNAL Prob_3_15_sva_2 : STD_LOGIC;
  SIGNAL Prob_6_14_1_sva_2 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL Prob_6_0_sva_2 : STD_LOGIC;
  SIGNAL Prob_6_15_sva_2 : STD_LOGIC;
  SIGNAL Prob_2_14_1_sva_2 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL Prob_2_0_sva_2 : STD_LOGIC;
  SIGNAL Prob_2_15_sva_2 : STD_LOGIC;
  SIGNAL Prob_7_14_1_sva_2 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL Prob_7_0_sva_2 : STD_LOGIC;
  SIGNAL Prob_7_15_sva_2 : STD_LOGIC;
  SIGNAL Prob_1_14_1_sva_2 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL Prob_1_0_sva_2 : STD_LOGIC;
  SIGNAL Prob_1_15_sva_2 : STD_LOGIC;
  SIGNAL Prob_8_14_1_sva_2 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL Prob_8_0_sva_2 : STD_LOGIC;
  SIGNAL Prob_8_15_sva_2 : STD_LOGIC;
  SIGNAL Prob_9_14_1_sva_2 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL Prob_9_0_sva_2 : STD_LOGIC;
  SIGNAL Prob_9_15_sva_2 : STD_LOGIC;
  SIGNAL perceptron_simple_k_7_0_sva_1 : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL k_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL FOR_B_lor_2_lpi_7_dfm_st : STD_LOGIC;
  SIGNAL FOR_B_2_lor_2_lpi_7_dfm_st : STD_LOGIC;
  SIGNAL FOR_B_4_lor_2_lpi_7_dfm_st : STD_LOGIC;
  SIGNAL CR1_simple_l_1_6_0_sva_5_0 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL CR2_simple_l_1_5_0_sva_4_0 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL Prob_0_sva_1_15 : STD_LOGIC;
  SIGNAL Prob_0_sva_1_14_1 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL Prob_0_sva_1_0 : STD_LOGIC;
  SIGNAL Prob_0_sva_2_15 : STD_LOGIC;
  SIGNAL Prob_0_sva_2_14_1 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL Prob_0_sva_2_0 : STD_LOGIC;
  SIGNAL MP3_simple_j_N_1_0_sva_1_1 : STD_LOGIC;
  SIGNAL MP3_simple_j_N_1_0_sva_0 : STD_LOGIC;
  SIGNAL MP3_simple_i_N_1_0_sva_1_1 : STD_LOGIC;
  SIGNAL MP3_simple_i_N_1_0_sva_0 : STD_LOGIC;
  SIGNAL CR1_simple_aux_15_lpi_7_mx1 : STD_LOGIC;
  SIGNAL CR1_simple_aux_14_1_lpi_7_mx1 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL CR1_simple_aux_0_lpi_7_mx1 : STD_LOGIC;
  SIGNAL FOR_B_acc_1_psp_sva_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL FOR_B_if_nor_ovfl_sva_1 : STD_LOGIC;
  SIGNAL FOR_B_if_and_unfl_sva_1 : STD_LOGIC;
  SIGNAL MP1_simple_bigger_lpi_6_mx1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL CR2_simple_aux_15_lpi_7_mx1 : STD_LOGIC;
  SIGNAL CR2_simple_aux_14_1_lpi_7_mx1 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL CR2_simple_aux_0_lpi_7_mx1 : STD_LOGIC;
  SIGNAL FOR_B_2_acc_1_psp_sva_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL FOR_B_2_if_nor_ovfl_sva_1 : STD_LOGIC;
  SIGNAL FOR_B_2_if_and_unfl_sva_1 : STD_LOGIC;
  SIGNAL MP2_simple_bigger_lpi_6_mx1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL CR3_simple_aux_15_lpi_7_mx1 : STD_LOGIC;
  SIGNAL CR3_simple_aux_14_1_lpi_7_mx1 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL CR3_simple_aux_0_lpi_7_mx1 : STD_LOGIC;
  SIGNAL FOR_B_4_acc_1_psp_1_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL MP3_simple_bigger_lpi_6_mx1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reshape_simple_add_N_10_0_lpi_4_mx0c1 : STD_LOGIC;
  SIGNAL perceptron_simple_k_7_0_sva_2 : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL FOR_K_7_FOR_K_7_nor_2_psp_sva_1 : STD_LOGIC;
  SIGNAL FOR_K_7_FOR_K_7_nor_1_psp_sva_1 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL FOR_K_7_nor_ovfl_sva_1 : STD_LOGIC;
  SIGNAL FOR_K_7_and_unfl_sva_1 : STD_LOGIC;
  SIGNAL max_sva_14_1_mx1 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL FOR_B_oelse_2_acc_itm_13 : STD_LOGIC;
  SIGNAL FOR_B_2_oelse_2_acc_itm_14 : STD_LOGIC;
  SIGNAL FOR_A_1_if_mux1h_4_cse : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL FOR_J_7_or_29_rgt : STD_LOGIC;
  SIGNAL FOR_J_7_and_81_rgt : STD_LOGIC;
  SIGNAL FOR_J_7_or_2_rgt : STD_LOGIC;
  SIGNAL FOR_J_7_and_27_rgt : STD_LOGIC;
  SIGNAL FOR_J_7_or_26_rgt : STD_LOGIC;
  SIGNAL FOR_J_7_and_75_rgt : STD_LOGIC;
  SIGNAL FOR_J_7_or_23_rgt : STD_LOGIC;
  SIGNAL FOR_J_7_and_69_rgt : STD_LOGIC;
  SIGNAL FOR_J_7_or_20_rgt : STD_LOGIC;
  SIGNAL FOR_J_7_and_63_rgt : STD_LOGIC;
  SIGNAL FOR_J_7_or_17_rgt : STD_LOGIC;
  SIGNAL FOR_J_7_and_57_rgt : STD_LOGIC;
  SIGNAL FOR_J_7_or_14_rgt : STD_LOGIC;
  SIGNAL FOR_J_7_and_51_rgt : STD_LOGIC;
  SIGNAL FOR_J_7_or_11_rgt : STD_LOGIC;
  SIGNAL FOR_J_7_and_45_rgt : STD_LOGIC;
  SIGNAL FOR_J_7_or_8_rgt : STD_LOGIC;
  SIGNAL FOR_J_7_and_39_rgt : STD_LOGIC;
  SIGNAL FOR_J_7_or_5_rgt : STD_LOGIC;
  SIGNAL FOR_J_7_and_33_rgt : STD_LOGIC;
  SIGNAL nand_cse_1 : STD_LOGIC;
  SIGNAL reg_FOR_I_asn_CR1_simple_add_AF_10_FOR_I_acc_psp_cse : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL reg_INIT_I_slc_INIT_I_acc_2_cse : STD_LOGIC;
  SIGNAL reg_FOR_I_2_acc_11_psp_cse : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL reg_FOR_I_2_acc_9_sdt_cse : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL reg_FOR_I_2_acc_10_psp_cse : STD_LOGIC;
  SIGNAL reg_FOR_I_2_acc_8_sdt_cse : STD_LOGIC;
  SIGNAL reg_FOR_I_4_acc_11_psp_cse : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL reg_FOR_I_4_acc_9_sdt_cse : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL reg_FOR_I_4_acc_8_sdt_2_0_cse : STD_LOGIC;
  SIGNAL FOR_I_nor_2_cse : STD_LOGIC;
  SIGNAL FOR_I_and_4_cse : STD_LOGIC;
  SIGNAL FOR_I_6_FOR_I_6_xnor_cse : STD_LOGIC;
  SIGNAL memory_1_or_2_cse : STD_LOGIC;
  SIGNAL memory_1_or_5_cse : STD_LOGIC;
  SIGNAL reg_FOR_A_1_lor_lpi_6_dfm_cse : STD_LOGIC;
  SIGNAL FOR_B_2_if_FOR_B_2_if_nor_cse : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL FOR_B_2_if_FOR_B_2_if_nor_1_cse : STD_LOGIC;
  SIGNAL memory_1_or_3_cse : STD_LOGIC;
  SIGNAL memory_1_or_12_cse : STD_LOGIC;
  SIGNAL memory_1_or_13_cse : STD_LOGIC;
  SIGNAL memory_1_or_6_cse_1 : STD_LOGIC;
  SIGNAL reshape_simple_add_N_or_cse : STD_LOGIC;
  SIGNAL reshape_simple_add_N_or_11_cse : STD_LOGIC;
  SIGNAL reshape_simple_add_N_or_2_cse : STD_LOGIC;
  SIGNAL FOR_I_nor_3_cse : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL FOR_I_nor_4_cse : STD_LOGIC;
  SIGNAL memory_1_or_17_cse : STD_LOGIC;
  SIGNAL memory_1_or_19_cse : STD_LOGIC;
  SIGNAL or_141_cse : STD_LOGIC;
  SIGNAL INIT_I_or_4_cse : STD_LOGIC;
  SIGNAL INIT_I_or_6_cse : STD_LOGIC;
  SIGNAL z_out_1_2 : STD_LOGIC;
  SIGNAL z_out_14_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL z_out_15_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL z_out_18_31_12 : STD_LOGIC_VECTOR (19 DOWNTO 0);
  SIGNAL z_out_27_2_0 : STD_LOGIC_VECTOR (2 DOWNTO 0);

  SIGNAL FOR_K_7_mux_1_nl : STD_LOGIC;
  SIGNAL FOR_K_7_mux_2_nl : STD_LOGIC;
  SIGNAL Prob_Prob_nor_nl : STD_LOGIC;
  SIGNAL Prob_and_19_nl : STD_LOGIC;
  SIGNAL FOR_K_7_mux_4_nl : STD_LOGIC;
  SIGNAL FOR_K_7_mux_5_nl : STD_LOGIC;
  SIGNAL Prob_Prob_nor_1_nl : STD_LOGIC;
  SIGNAL Prob_and_17_nl : STD_LOGIC;
  SIGNAL FOR_K_7_mux_7_nl : STD_LOGIC;
  SIGNAL FOR_K_7_mux_8_nl : STD_LOGIC;
  SIGNAL Prob_Prob_nor_2_nl : STD_LOGIC;
  SIGNAL Prob_and_15_nl : STD_LOGIC;
  SIGNAL FOR_K_7_mux_10_nl : STD_LOGIC;
  SIGNAL FOR_K_7_mux_11_nl : STD_LOGIC;
  SIGNAL Prob_Prob_nor_3_nl : STD_LOGIC;
  SIGNAL Prob_and_13_nl : STD_LOGIC;
  SIGNAL FOR_K_7_mux_13_nl : STD_LOGIC;
  SIGNAL FOR_K_7_mux_14_nl : STD_LOGIC;
  SIGNAL Prob_Prob_nor_4_nl : STD_LOGIC;
  SIGNAL Prob_and_11_nl : STD_LOGIC;
  SIGNAL FOR_K_7_mux_16_nl : STD_LOGIC;
  SIGNAL FOR_K_7_mux_17_nl : STD_LOGIC;
  SIGNAL Prob_Prob_nor_5_nl : STD_LOGIC;
  SIGNAL Prob_and_9_nl : STD_LOGIC;
  SIGNAL FOR_K_7_mux_19_nl : STD_LOGIC;
  SIGNAL FOR_K_7_mux_20_nl : STD_LOGIC;
  SIGNAL Prob_Prob_nor_6_nl : STD_LOGIC;
  SIGNAL Prob_and_7_nl : STD_LOGIC;
  SIGNAL FOR_K_7_mux_22_nl : STD_LOGIC;
  SIGNAL FOR_K_7_mux_23_nl : STD_LOGIC;
  SIGNAL Prob_Prob_nor_7_nl : STD_LOGIC;
  SIGNAL Prob_and_5_nl : STD_LOGIC;
  SIGNAL FOR_K_7_mux_25_nl : STD_LOGIC;
  SIGNAL FOR_K_7_mux_26_nl : STD_LOGIC;
  SIGNAL Prob_Prob_nor_8_nl : STD_LOGIC;
  SIGNAL Prob_and_3_nl : STD_LOGIC;
  SIGNAL CR1_simple_l_not_1_nl : STD_LOGIC;
  SIGNAL CR1_simple_j_not_nl : STD_LOGIC;
  SIGNAL CR1_simple_i_nor_nl : STD_LOGIC;
  SIGNAL CR1_simple_aux_mux_14_nl : STD_LOGIC;
  SIGNAL CR1_simple_aux_mux_13_nl : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL not_410_nl : STD_LOGIC;
  SIGNAL CR1_simple_aux_mux_12_nl : STD_LOGIC;
  SIGNAL not_408_nl : STD_LOGIC;
  SIGNAL MP1_simple_i_not_nl : STD_LOGIC;
  SIGNAL MP1_simple_i_N_not_nl : STD_LOGIC;
  SIGNAL MP1_simple_a_nor_nl : STD_LOGIC;
  SIGNAL MP1_simple_b_not_nl : STD_LOGIC;
  SIGNAL memory_1_mux_3_nl : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL MP1_simple_bigger_not_nl : STD_LOGIC;
  SIGNAL CR1_simple_aux_mux_11_nl : STD_LOGIC;
  SIGNAL CR1_simple_aux_mux_10_nl : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL not_406_nl : STD_LOGIC;
  SIGNAL CR1_simple_aux_mux_9_nl : STD_LOGIC;
  SIGNAL not_404_nl : STD_LOGIC;
  SIGNAL MP2_simple_i_not_nl : STD_LOGIC;
  SIGNAL MP2_simple_i_N_not_nl : STD_LOGIC;
  SIGNAL MP2_simple_a_nor_nl : STD_LOGIC;
  SIGNAL MP2_simple_b_not_nl : STD_LOGIC;
  SIGNAL memory_1_mux_4_nl : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL MP2_simple_bigger_not_nl : STD_LOGIC;
  SIGNAL CR1_simple_aux_mux_8_nl : STD_LOGIC;
  SIGNAL CR1_simple_aux_mux_7_nl : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL not_402_nl : STD_LOGIC;
  SIGNAL CR1_simple_aux_mux_6_nl : STD_LOGIC;
  SIGNAL MP3_simple_i_not_nl : STD_LOGIC;
  SIGNAL MP3_simple_a_not_nl : STD_LOGIC;
  SIGNAL MP3_simple_b_not_nl : STD_LOGIC;
  SIGNAL memory_1_mux_5_nl : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL MP3_simple_bigger_not_nl : STD_LOGIC;
  SIGNAL FOR_K_7_mux_28_nl : STD_LOGIC;
  SIGNAL FOR_K_7_mux_29_nl : STD_LOGIC;
  SIGNAL Prob_Prob_nor_9_nl : STD_LOGIC;
  SIGNAL Prob_and_1_nl : STD_LOGIC;
  SIGNAL FOR_K_7_acc_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL for_mux_1_nl : STD_LOGIC;
  SIGNAL for_mux_2_nl : STD_LOGIC;
  SIGNAL FOR_B_if_FOR_B_if_nor_nl : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL FOR_B_if_nor_2_nl : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL FOR_B_if_FOR_B_if_nor_1_nl : STD_LOGIC;
  SIGNAL FOR_B_oelse_2_acc_nl : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL FOR_B_oelse_acc_nl : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL FOR_B_2_if_nor_2_nl : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL FOR_B_2_oelse_2_acc_nl : STD_LOGIC_VECTOR (14 DOWNTO 0);
  SIGNAL FOR_B_2_oelse_acc_nl : STD_LOGIC_VECTOR (14 DOWNTO 0);
  SIGNAL FOR_B_4_if_acc_12_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL FOR_B_4_if_acc_9_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL FOR_B_4_oelse_acc_nl : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL FOR_K_7_nor_3_nl : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL BIAS_I_BIAS_I_and_2_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL FOR_B_if_asn_CR1_simple_add_M_10_FOR_B_if_acc_nl : STD_LOGIC_VECTOR (4 DOWNTO
      0);
  SIGNAL FOR_K_FOR_K_and_5_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL BIAS_I_BIAS_I_and_3_nl : STD_LOGIC;
  SIGNAL BIAS_I_2_BIAS_I_2_and_3_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL FOR_K_FOR_K_and_4_nl : STD_LOGIC;
  SIGNAL FOR_K_FOR_K_and_11_nl : STD_LOGIC;
  SIGNAL BIAS_I_2_BIAS_I_2_and_2_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL CR1_simple_l_CR1_simple_l_and_1_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL CR1_simple_l_nor_nl : STD_LOGIC;
  SIGNAL B_1_nor_nl : STD_LOGIC;
  SIGNAL BIAS_I_2_BIAS_I_2_and_1_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL BIAS_I_BIAS_I_and_1_nl : STD_LOGIC;
  SIGNAL CR2_simple_k_CR2_simple_k_and_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL CR2_simple_k_not_nl : STD_LOGIC;
  SIGNAL CR2_simple_l_CR2_simple_l_and_1_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL CR2_simple_l_not_nl : STD_LOGIC;
  SIGNAL B_2_nor_nl : STD_LOGIC;
  SIGNAL FOR_K_FOR_K_and_3_nl : STD_LOGIC;
  SIGNAL FOR_K_FOR_K_and_10_nl : STD_LOGIC;
  SIGNAL BIAS_I_1_BIAS_I_1_and_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL BIAS_I_2_BIAS_I_2_and_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL FOR_K_FOR_K_and_2_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL FOR_K_FOR_K_and_1_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL B_3_nor_nl : STD_LOGIC;
  SIGNAL FOR_K_7_FOR_K_7_and_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL FOR_K_7_acc_9_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL FOR_K_FOR_K_and_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL BIAS_I_BIAS_I_and_nl : STD_LOGIC;
  SIGNAL memory_1_and_1_nl : STD_LOGIC;
  SIGNAL memory_1_mux1h_1_nl : STD_LOGIC;
  SIGNAL memory_1_and_4_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL memory_1_mux1h_5_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL memory_1_mux1h_12_nl : STD_LOGIC;
  SIGNAL memory_1_mux1h_13_nl : STD_LOGIC;
  SIGNAL memory_1_and_5_nl : STD_LOGIC;
  SIGNAL memory_1_mux1h_6_nl : STD_LOGIC;
  SIGNAL memory_1_and_6_nl : STD_LOGIC;
  SIGNAL memory_1_mux1h_7_nl : STD_LOGIC;
  SIGNAL memory_1_and_7_nl : STD_LOGIC;
  SIGNAL memory_1_mux1h_8_nl : STD_LOGIC;
  SIGNAL memory_1_and_8_nl : STD_LOGIC;
  SIGNAL memory_1_mux1h_9_nl : STD_LOGIC;
  SIGNAL reshape_simple_add_N_and_nl : STD_LOGIC;
  SIGNAL reshape_simple_add_N_mux1h_nl : STD_LOGIC;
  SIGNAL reshape_simple_add_N_and_2_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL reshape_simple_add_N_mux1h_4_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL reshape_simple_add_N_mux1h_9_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL reshape_simple_add_N_or_3_nl : STD_LOGIC;
  SIGNAL reshape_simple_add_N_or_15_nl : STD_LOGIC;
  SIGNAL reshape_simple_add_N_and_3_nl : STD_LOGIC;
  SIGNAL reshape_simple_add_N_mux1h_5_nl : STD_LOGIC;
  SIGNAL reshape_simple_add_N_and_4_nl : STD_LOGIC;
  SIGNAL reshape_simple_add_N_mux1h_6_nl : STD_LOGIC;
  SIGNAL reshape_simple_add_N_and_5_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL reshape_simple_add_N_mux1h_7_nl : STD_LOGIC;
  SIGNAL reshape_simple_add_N_mux1h_10_nl : STD_LOGIC;
  SIGNAL memory_1_and_nl : STD_LOGIC;
  SIGNAL memory_1_memory_1_mux_nl : STD_LOGIC;
  SIGNAL memory_1_and_9_nl : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL memory_1_mux1h_10_nl : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL FOR_I_FOR_I_nor_1_nl : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL BIAS_I_BIAS_I_nor_nl : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL memory_1_and_10_nl : STD_LOGIC;
  SIGNAL memory_1_mux1h_11_nl : STD_LOGIC;
  SIGNAL FOR_I_FOR_I_nor_2_nl : STD_LOGIC;
  SIGNAL BIAS_I_BIAS_I_nor_3_nl : STD_LOGIC;
  SIGNAL memory_2_and_3_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL memory_2_mux1h_1_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL FOR_B_2_if_acc_12_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL FOR_B_4_if_acc_16_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL memory_2_not_4_nl : STD_LOGIC;
  SIGNAL memory_2_and_4_nl : STD_LOGIC;
  SIGNAL memory_2_mux1h_4_nl : STD_LOGIC;
  SIGNAL memory_2_and_5_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL memory_2_mux1h_5_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL memory_2_not_6_nl : STD_LOGIC;
  SIGNAL memory_2_and_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL memory_2_mux1h_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL FOR_B_1_if_acc_5_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL FOR_B_3_if_acc_5_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL memory_2_not_1_nl : STD_LOGIC;
  SIGNAL memory_2_and_1_nl : STD_LOGIC;
  SIGNAL memory_2_mux1h_2_nl : STD_LOGIC;
  SIGNAL memory_2_and_2_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL memory_2_mux1h_3_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL memory_2_not_3_nl : STD_LOGIC;
  SIGNAL MP1_simple_bigger_mux1h_nl : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL or_198_nl : STD_LOGIC;
  SIGNAL memory_2_nand_nl : STD_LOGIC;
  SIGNAL acc_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL INIT_I_mux1h_7_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL INIT_I_or_13_nl : STD_LOGIC;
  SIGNAL INIT_I_or_14_nl : STD_LOGIC;
  SIGNAL INIT_I_or_15_nl : STD_LOGIC;
  SIGNAL INIT_I_nor_1_nl : STD_LOGIC;
  SIGNAL INIT_I_mux1h_8_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL INIT_I_or_17_nl : STD_LOGIC;
  SIGNAL acc_1_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL FOR_A_1_if_mux1h_9_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL FOR_A_3_if_acc_16_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL FOR_A_1_if_nor_3_nl : STD_LOGIC;
  SIGNAL FOR_A_1_if_FOR_A_1_if_or_1_nl : STD_LOGIC;
  SIGNAL FOR_B_mux1h_6_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL FOR_B_or_3_nl : STD_LOGIC;
  SIGNAL FOR_B_FOR_B_mux_1_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL FOR_B_if_mux1h_6_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL FOR_B_if_or_4_nl : STD_LOGIC;
  SIGNAL FOR_B_if_mux1h_7_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL acc_4_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL FOR_A_1_if_mux1h_10_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL FOR_A_1_if_and_1_nl : STD_LOGIC;
  SIGNAL FOR_A_1_if_mux1h_11_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL FOR_J_1_mux1h_2_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL FOR_J_3_mux1h_2_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL FOR_K_6_mux1h_2_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL FOR_K_6_or_5_nl : STD_LOGIC;
  SIGNAL mux1h_1_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL or_nl : STD_LOGIC;
  SIGNAL or_663_nl : STD_LOGIC;
  SIGNAL FOR_A_1_if_FOR_A_1_if_and_1_nl : STD_LOGIC;
  SIGNAL FOR_A_1_if_mux1h_12_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL INIT_J_mux1h_2_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL INIT_I_mux1h_9_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL INIT_I_or_18_nl : STD_LOGIC;
  SIGNAL INIT_I_mux1h_10_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL FOR_A_3_if_acc_17_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL INIT_I_or_19_nl : STD_LOGIC;
  SIGNAL FOR_B_4_if_mux_2_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL FOR_B_4_if_mux_3_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL INIT_I_mux1h_11_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL INIT_I_mux1h_12_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL INIT_L_mux1h_2_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL FOR_B_mux1h_7_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL FOR_B_mux1h_8_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL FOR_B_mux1h_9_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL FOR_B_mux1h_10_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL FOR_B_or_4_nl : STD_LOGIC;
  SIGNAL FOR_B_if_mux1h_8_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL FOR_B_if_mux1h_9_nl : STD_LOGIC;
  SIGNAL mul_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL FOR_B_if_mux1h_10_nl : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL FOR_B_if_mux1h_11_nl : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL FOR_B_if_or_5_nl : STD_LOGIC;
  SIGNAL FOR_A_5_if_mux_1_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL acc_21_nl : STD_LOGIC_VECTOR (17 DOWNTO 0);
  SIGNAL FOR_I_mux1h_2_nl : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL FOR_I_or_3_nl : STD_LOGIC;
  SIGNAL FOR_I_nor_5_nl : STD_LOGIC;
  SIGNAL FOR_I_mux1h_3_nl : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL FOR_I_or_5_nl : STD_LOGIC;
  SIGNAL FOR_B_2_if_mux_4_nl : STD_LOGIC;
  SIGNAL FOR_B_2_if_mux_5_nl : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL FOR_B_2_if_mux_6_nl : STD_LOGIC;
  SIGNAL FOR_A_3_if_mux_2_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL FOR_A_5_if_acc_21_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL FOR_A_3_if_mux_3_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL FOR_B_3_if_mux1h_2_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL FOR_B_3_if_FOR_B_3_if_mux_1_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL FOR_B_3_if_or_1_nl : STD_LOGIC;
  SIGNAL INIT_I_2_mux1h_2_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL INIT_I_2_mux1h_3_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL index_rsci_idat_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL index_rsci_dat : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT CNN_main_simple_core_core_fsm
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      fsm_output : OUT STD_LOGIC_VECTOR (91 DOWNTO 0);
      INIT_I_C_1_tr0 : IN STD_LOGIC;
      INIT_J_C_0_tr0 : IN STD_LOGIC;
      INIT_L_C_0_tr0 : IN STD_LOGIC;
      FOR_B_C_1_tr0 : IN STD_LOGIC;
      FOR_A_C_0_tr0 : IN STD_LOGIC;
      FOR_I_C_2_tr0 : IN STD_LOGIC;
      FOR_J_C_0_tr0 : IN STD_LOGIC;
      FOR_K_C_0_tr0 : IN STD_LOGIC;
      BIAS_I_C_2_tr0 : IN STD_LOGIC;
      BIAS_J_C_0_tr0 : IN STD_LOGIC;
      FOR_L_C_0_tr0 : IN STD_LOGIC;
      FOR_A_1_C_1_tr0 : IN STD_LOGIC;
      FOR_B_1_C_1_tr0 : IN STD_LOGIC;
      FOR_I_1_C_1_tr0 : IN STD_LOGIC;
      FOR_J_1_C_1_tr0 : IN STD_LOGIC;
      FOR_K_1_C_0_tr0 : IN STD_LOGIC;
      INIT_I_1_C_1_tr0 : IN STD_LOGIC;
      INIT_J_1_C_0_tr0 : IN STD_LOGIC;
      INIT_L_1_C_0_tr0 : IN STD_LOGIC;
      FOR_B_2_C_1_tr0 : IN STD_LOGIC;
      FOR_A_2_C_0_tr0 : IN STD_LOGIC;
      FOR_I_2_C_2_tr0 : IN STD_LOGIC;
      FOR_J_2_C_0_tr0 : IN STD_LOGIC;
      FOR_K_2_C_0_tr0 : IN STD_LOGIC;
      BIAS_I_1_C_2_tr0 : IN STD_LOGIC;
      BIAS_J_1_C_0_tr0 : IN STD_LOGIC;
      FOR_L_1_C_0_tr0 : IN STD_LOGIC;
      FOR_A_3_C_1_tr0 : IN STD_LOGIC;
      FOR_B_3_C_1_tr0 : IN STD_LOGIC;
      FOR_I_3_C_1_tr0 : IN STD_LOGIC;
      FOR_J_3_C_1_tr0 : IN STD_LOGIC;
      FOR_K_3_C_0_tr0 : IN STD_LOGIC;
      INIT_I_2_C_1_tr0 : IN STD_LOGIC;
      INIT_J_2_C_0_tr0 : IN STD_LOGIC;
      INIT_L_2_C_0_tr0 : IN STD_LOGIC;
      FOR_B_4_C_1_tr0 : IN STD_LOGIC;
      FOR_A_4_C_0_tr0 : IN STD_LOGIC;
      FOR_I_4_C_2_tr0 : IN STD_LOGIC;
      FOR_J_4_C_0_tr0 : IN STD_LOGIC;
      FOR_K_4_C_0_tr0 : IN STD_LOGIC;
      BIAS_I_2_C_2_tr0 : IN STD_LOGIC;
      BIAS_J_2_C_0_tr0 : IN STD_LOGIC;
      FOR_L_2_C_0_tr0 : IN STD_LOGIC;
      FOR_A_5_C_1_tr0 : IN STD_LOGIC;
      FOR_B_5_C_1_tr0 : IN STD_LOGIC;
      FOR_I_5_C_1_tr0 : IN STD_LOGIC;
      FOR_J_5_C_1_tr0 : IN STD_LOGIC;
      FOR_K_5_C_0_tr0 : IN STD_LOGIC;
      FOR_K_6_C_2_tr0 : IN STD_LOGIC;
      FOR_J_6_C_0_tr0 : IN STD_LOGIC;
      FOR_I_6_C_0_tr0 : IN STD_LOGIC;
      FOR_K_7_C_1_tr0 : IN STD_LOGIC;
      FOR_J_7_C_1_tr0 : IN STD_LOGIC;
      for_C_0_tr0 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL CNN_main_simple_core_core_fsm_inst_fsm_output : STD_LOGIC_VECTOR (91 DOWNTO
      0);
  SIGNAL CNN_main_simple_core_core_fsm_inst_INIT_I_C_1_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_INIT_J_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_INIT_L_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_B_C_1_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_A_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_I_C_2_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_J_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_BIAS_I_C_2_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_BIAS_J_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_L_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_A_1_C_1_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_B_1_C_1_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_I_1_C_1_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_J_1_C_1_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_K_1_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_INIT_I_1_C_1_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_INIT_J_1_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_INIT_L_1_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_B_2_C_1_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_A_2_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_I_2_C_2_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_J_2_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_K_2_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_BIAS_I_1_C_2_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_BIAS_J_1_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_L_1_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_A_3_C_1_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_B_3_C_1_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_I_3_C_1_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_J_3_C_1_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_K_3_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_INIT_I_2_C_1_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_INIT_J_2_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_INIT_L_2_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_B_4_C_1_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_A_4_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_I_4_C_2_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_J_4_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_K_4_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_BIAS_I_2_C_2_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_BIAS_J_2_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_L_2_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_A_5_C_1_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_B_5_C_1_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_I_5_C_1_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_J_5_C_1_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_K_5_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_K_6_C_2_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_J_6_C_0_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_K_7_C_1_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_FOR_J_7_C_1_tr0 : STD_LOGIC;
  SIGNAL CNN_main_simple_core_core_fsm_inst_for_C_0_tr0 : STD_LOGIC;

  FUNCTION CONV_SL_1_1(input:BOOLEAN)
  RETURN STD_LOGIC IS
  BEGIN
    IF input THEN RETURN '1';ELSE RETURN '0';END IF;
  END;

  FUNCTION MUX1HOT_s_1_10_2(input_9 : STD_LOGIC;
  input_8 : STD_LOGIC;
  input_7 : STD_LOGIC;
  input_6 : STD_LOGIC;
  input_5 : STD_LOGIC;
  input_4 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(9 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
      tmp := sel(4);
      result := result or ( input_4 and tmp);
      tmp := sel(5);
      result := result or ( input_5 and tmp);
      tmp := sel(6);
      result := result or ( input_6 and tmp);
      tmp := sel(7);
      result := result or ( input_7 and tmp);
      tmp := sel(8);
      result := result or ( input_8 and tmp);
      tmp := sel(9);
      result := result or ( input_9 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_3_2(input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_4_2(input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_5_2(input_4 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
      tmp := sel(4);
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_7_2(input_6 : STD_LOGIC;
  input_5 : STD_LOGIC;
  input_4 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(6 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
      tmp := sel(4);
      result := result or ( input_4 and tmp);
      tmp := sel(5);
      result := result or ( input_5 and tmp);
      tmp := sel(6);
      result := result or ( input_6 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_8_2(input_7 : STD_LOGIC;
  input_6 : STD_LOGIC;
  input_5 : STD_LOGIC;
  input_4 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(7 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
      tmp := sel(4);
      result := result or ( input_4 and tmp);
      tmp := sel(5);
      result := result or ( input_5 and tmp);
      tmp := sel(6);
      result := result or ( input_6 and tmp);
      tmp := sel(7);
      result := result or ( input_7 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_9_2(input_8 : STD_LOGIC;
  input_7 : STD_LOGIC;
  input_6 : STD_LOGIC;
  input_5 : STD_LOGIC;
  input_4 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(8 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
      tmp := sel(4);
      result := result or ( input_4 and tmp);
      tmp := sel(5);
      result := result or ( input_5 and tmp);
      tmp := sel(6);
      result := result or ( input_6 and tmp);
      tmp := sel(7);
      result := result or ( input_7 and tmp);
      tmp := sel(8);
      result := result or ( input_8 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_14_3_2(input_2 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(13 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(13 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_16_3_2(input_2 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(15 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(15 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_16_4_2(input_3 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(15 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(15 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_16_6_2(input_5 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(15 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(15 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_16_9_2(input_8 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(8 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(15 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(15 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_2_19_2(input_18 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_17 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(18 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(1 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(1 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
      tmp := (OTHERS=>sel( 17));
      result := result or ( input_17 and tmp);
      tmp := (OTHERS=>sel( 18));
      result := result or ( input_18 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_2_3_2(input_2 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(1 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(1 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_2_4_2(input_3 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(1 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(1 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_2_5_2(input_4 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(1 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(1 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_2_7_2(input_6 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(6 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(1 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(1 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_3_10_2(input_9 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(9 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_3_3_2(input_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_3_4_2(input_3 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_3_5_2(input_4 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_4_12_2(input_11 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(11 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_4_5_2(input_4 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_4_6_2(input_5 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_4_7_2(input_6 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(6 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_5_10_2(input_9 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(9 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_5_6_2(input_5 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_5_7_2(input_6 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(6 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_6_4_2(input_3 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_8_3_2(input_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(7 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(7 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX_s_1_10_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_4 : STD_LOGIC;
  input_5 : STD_LOGIC;
  input_6 : STD_LOGIC;
  input_7 : STD_LOGIC;
  input_8 : STD_LOGIC;
  input_9 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN "0000" =>
          result := input_0;
        WHEN "0001" =>
          result := input_1;
        WHEN "0010" =>
          result := input_2;
        WHEN "0011" =>
          result := input_3;
        WHEN "0100" =>
          result := input_4;
        WHEN "0101" =>
          result := input_5;
        WHEN "0110" =>
          result := input_6;
        WHEN "0111" =>
          result := input_7;
        WHEN "1000" =>
          result := input_8;
        WHEN others =>
          result := input_9;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_s_1_2_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  sel : STD_LOGIC)
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_11_2_2(input_0 : STD_LOGIC_VECTOR(10 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(10 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(10 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(10 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_14_10_2(input_0 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(13 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(13 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN "0000" =>
          result := input_0;
        WHEN "0001" =>
          result := input_1;
        WHEN "0010" =>
          result := input_2;
        WHEN "0011" =>
          result := input_3;
        WHEN "0100" =>
          result := input_4;
        WHEN "0101" =>
          result := input_5;
        WHEN "0110" =>
          result := input_6;
        WHEN "0111" =>
          result := input_7;
        WHEN "1000" =>
          result := input_8;
        WHEN others =>
          result := input_9;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_14_2_2(input_0 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(13 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(13 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(13 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_16_2_2(input_0 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(15 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(15 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_2_2_2(input_0 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(1 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(1 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_3_2_2(input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_4_2_2(input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_6_2_2(input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_8_2_2(input_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(7 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(7 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION READSLICE_17_18(input:STD_LOGIC_VECTOR(17 DOWNTO 0);index:INTEGER)
  RETURN STD_LOGIC_VECTOR IS
    CONSTANT slice_exes:STD_LOGIC_VECTOR(16 DOWNTO 0):=(OTHERS=>'X');
    CONSTANT left_range:INTEGER:=index+16;
  BEGIN
    IF index<0 OR 1<index THEN
      RETURN slice_exes;
    END IF;
    RETURN input(left_range DOWNTO index);
  END;

  FUNCTION READSLICE_1_14(input:STD_LOGIC_VECTOR(13 DOWNTO 0);index:INTEGER)
  RETURN STD_LOGIC IS
  BEGIN
    IF index<0 OR 13<index THEN
      RETURN 'X';
    END IF;
    RETURN input(index);
  END;

  FUNCTION READSLICE_1_15(input:STD_LOGIC_VECTOR(14 DOWNTO 0);index:INTEGER)
  RETURN STD_LOGIC IS
  BEGIN
    IF index<0 OR 14<index THEN
      RETURN 'X';
    END IF;
    RETURN input(index);
  END;

  FUNCTION READSLICE_1_16(input:STD_LOGIC_VECTOR(15 DOWNTO 0);index:INTEGER)
  RETURN STD_LOGIC IS
  BEGIN
    IF index<0 OR 15<index THEN
      RETURN 'X';
    END IF;
    RETURN input(index);
  END;

  FUNCTION READSLICE_1_4(input:STD_LOGIC_VECTOR(3 DOWNTO 0);index:INTEGER)
  RETURN STD_LOGIC IS
  BEGIN
    IF index<0 OR 3<index THEN
      RETURN 'X';
    END IF;
    RETURN input(index);
  END;

  FUNCTION READSLICE_1_7(input:STD_LOGIC_VECTOR(6 DOWNTO 0);index:INTEGER)
  RETURN STD_LOGIC IS
  BEGIN
    IF index<0 OR 6<index THEN
      RETURN 'X';
    END IF;
    RETURN input(index);
  END;

  FUNCTION READSLICE_20_32(input:STD_LOGIC_VECTOR(31 DOWNTO 0);index:INTEGER)
  RETURN STD_LOGIC_VECTOR IS
    CONSTANT slice_exes:STD_LOGIC_VECTOR(19 DOWNTO 0):=(OTHERS=>'X');
    CONSTANT left_range:INTEGER:=index+19;
  BEGIN
    IF index<0 OR 12<index THEN
      RETURN slice_exes;
    END IF;
    RETURN input(left_range DOWNTO index);
  END;

  FUNCTION READSLICE_2_3(input:STD_LOGIC_VECTOR(2 DOWNTO 0);index:INTEGER)
  RETURN STD_LOGIC_VECTOR IS
    CONSTANT slice_exes:STD_LOGIC_VECTOR(1 DOWNTO 0):=(OTHERS=>'X');
    CONSTANT left_range:INTEGER:=index+1;
  BEGIN
    IF index<0 OR 1<index THEN
      RETURN slice_exes;
    END IF;
    RETURN input(left_range DOWNTO index);
  END;

  FUNCTION READSLICE_3_4(input:STD_LOGIC_VECTOR(3 DOWNTO 0);index:INTEGER)
  RETURN STD_LOGIC_VECTOR IS
    CONSTANT slice_exes:STD_LOGIC_VECTOR(2 DOWNTO 0):=(OTHERS=>'X');
    CONSTANT left_range:INTEGER:=index+2;
  BEGIN
    IF index<0 OR 1<index THEN
      RETURN slice_exes;
    END IF;
    RETURN input(left_range DOWNTO index);
  END;

BEGIN
  -- Default Constant Signal Assignments

  index_rsci : work.ccs_out_pkg_v1.ccs_out_v1
    GENERIC MAP(
      rscid => 10,
      width => 4
      )
    PORT MAP(
      idat => index_rsci_idat_1,
      dat => index_rsci_dat
    );
  index_rsci_idat_1 <= index_rsci_idat;
  index_rsc_dat <= index_rsci_dat;

  image_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_index_rsc_triosy_obj_ld_cse,
      lz => image_rsc_triosy_lz
    );
  F_1_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_index_rsc_triosy_obj_ld_cse,
      lz => F_1_rsc_triosy_lz
    );
  B_1_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_index_rsc_triosy_obj_ld_cse,
      lz => B_1_rsc_triosy_lz
    );
  F_2_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_index_rsc_triosy_obj_ld_cse,
      lz => F_2_rsc_triosy_lz
    );
  B_2_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_index_rsc_triosy_obj_ld_cse,
      lz => B_2_rsc_triosy_lz
    );
  F_3_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_index_rsc_triosy_obj_ld_cse,
      lz => F_3_rsc_triosy_lz
    );
  B_3_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_index_rsc_triosy_obj_ld_cse,
      lz => B_3_rsc_triosy_lz
    );
  P_W_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_index_rsc_triosy_obj_ld_cse,
      lz => P_W_rsc_triosy_lz
    );
  P_B_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_index_rsc_triosy_obj_ld_cse,
      lz => P_B_rsc_triosy_lz
    );
  index_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_index_rsc_triosy_obj_ld_cse,
      lz => index_rsc_triosy_lz
    );
  CNN_main_simple_core_core_fsm_inst : CNN_main_simple_core_core_fsm
    PORT MAP(
      clk => clk,
      rst => rst,
      fsm_output => CNN_main_simple_core_core_fsm_inst_fsm_output,
      INIT_I_C_1_tr0 => CNN_main_simple_core_core_fsm_inst_INIT_I_C_1_tr0,
      INIT_J_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_INIT_J_C_0_tr0,
      INIT_L_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_INIT_L_C_0_tr0,
      FOR_B_C_1_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_B_C_1_tr0,
      FOR_A_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_A_C_0_tr0,
      FOR_I_C_2_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_I_C_2_tr0,
      FOR_J_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_J_C_0_tr0,
      FOR_K_C_0_tr0 => FOR_I_6_FOR_I_6_xnor_cse,
      BIAS_I_C_2_tr0 => CNN_main_simple_core_core_fsm_inst_BIAS_I_C_2_tr0,
      BIAS_J_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_BIAS_J_C_0_tr0,
      FOR_L_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_L_C_0_tr0,
      FOR_A_1_C_1_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_A_1_C_1_tr0,
      FOR_B_1_C_1_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_B_1_C_1_tr0,
      FOR_I_1_C_1_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_I_1_C_1_tr0,
      FOR_J_1_C_1_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_J_1_C_1_tr0,
      FOR_K_1_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_K_1_C_0_tr0,
      INIT_I_1_C_1_tr0 => CNN_main_simple_core_core_fsm_inst_INIT_I_1_C_1_tr0,
      INIT_J_1_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_INIT_J_1_C_0_tr0,
      INIT_L_1_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_INIT_L_1_C_0_tr0,
      FOR_B_2_C_1_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_B_2_C_1_tr0,
      FOR_A_2_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_A_2_C_0_tr0,
      FOR_I_2_C_2_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_I_2_C_2_tr0,
      FOR_J_2_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_J_2_C_0_tr0,
      FOR_K_2_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_K_2_C_0_tr0,
      BIAS_I_1_C_2_tr0 => CNN_main_simple_core_core_fsm_inst_BIAS_I_1_C_2_tr0,
      BIAS_J_1_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_BIAS_J_1_C_0_tr0,
      FOR_L_1_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_L_1_C_0_tr0,
      FOR_A_3_C_1_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_A_3_C_1_tr0,
      FOR_B_3_C_1_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_B_3_C_1_tr0,
      FOR_I_3_C_1_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_I_3_C_1_tr0,
      FOR_J_3_C_1_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_J_3_C_1_tr0,
      FOR_K_3_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_K_3_C_0_tr0,
      INIT_I_2_C_1_tr0 => CNN_main_simple_core_core_fsm_inst_INIT_I_2_C_1_tr0,
      INIT_J_2_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_INIT_J_2_C_0_tr0,
      INIT_L_2_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_INIT_L_2_C_0_tr0,
      FOR_B_4_C_1_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_B_4_C_1_tr0,
      FOR_A_4_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_A_4_C_0_tr0,
      FOR_I_4_C_2_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_I_4_C_2_tr0,
      FOR_J_4_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_J_4_C_0_tr0,
      FOR_K_4_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_K_4_C_0_tr0,
      BIAS_I_2_C_2_tr0 => CNN_main_simple_core_core_fsm_inst_BIAS_I_2_C_2_tr0,
      BIAS_J_2_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_BIAS_J_2_C_0_tr0,
      FOR_L_2_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_L_2_C_0_tr0,
      FOR_A_5_C_1_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_A_5_C_1_tr0,
      FOR_B_5_C_1_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_B_5_C_1_tr0,
      FOR_I_5_C_1_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_I_5_C_1_tr0,
      FOR_J_5_C_1_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_J_5_C_1_tr0,
      FOR_K_5_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_K_5_C_0_tr0,
      FOR_K_6_C_2_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_K_6_C_2_tr0,
      FOR_J_6_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_J_6_C_0_tr0,
      FOR_I_6_C_0_tr0 => FOR_I_6_FOR_I_6_xnor_cse,
      FOR_K_7_C_1_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_K_7_C_1_tr0,
      FOR_J_7_C_1_tr0 => CNN_main_simple_core_core_fsm_inst_FOR_J_7_C_1_tr0,
      for_C_0_tr0 => CNN_main_simple_core_core_fsm_inst_for_C_0_tr0
    );
  fsm_output <= CNN_main_simple_core_core_fsm_inst_fsm_output;
  CNN_main_simple_core_core_fsm_inst_INIT_I_C_1_tr0 <= NOT reg_INIT_I_slc_INIT_I_acc_2_cse;
  CNN_main_simple_core_core_fsm_inst_INIT_J_C_0_tr0 <= NOT (z_out(2));
  CNN_main_simple_core_core_fsm_inst_INIT_L_C_0_tr0 <= z_out_13(6);
  CNN_main_simple_core_core_fsm_inst_FOR_B_C_1_tr0 <= NOT((CR1_simple_b_1_0_sva_1(0))
      XOR (CR1_simple_b_1_0_sva_1(1)));
  CNN_main_simple_core_core_fsm_inst_FOR_A_C_0_tr0 <= NOT((z_out_2(0)) XOR (z_out_2(1)));
  CNN_main_simple_core_core_fsm_inst_FOR_I_C_2_tr0 <= NOT FOR_I_slc_FOR_I_acc_2_itm;
  CNN_main_simple_core_core_fsm_inst_FOR_J_C_0_tr0 <= NOT (z_out(2));
  CNN_main_simple_core_core_fsm_inst_BIAS_I_C_2_tr0 <= NOT BIAS_I_slc_BIAS_I_acc_2_itm;
  CNN_main_simple_core_core_fsm_inst_BIAS_J_C_0_tr0 <= NOT (z_out(2));
  CNN_main_simple_core_core_fsm_inst_FOR_L_C_0_tr0 <= z_out_13(6);
  CNN_main_simple_core_core_fsm_inst_FOR_A_1_C_1_tr0 <= NOT((CR1_simple_b_1_0_sva_1(0))
      XOR (CR1_simple_b_1_0_sva_1(1)));
  CNN_main_simple_core_core_fsm_inst_FOR_B_1_C_1_tr0 <= NOT((CR1_simple_b_1_0_sva_1(0))
      XOR (CR1_simple_b_1_0_sva_1(1)));
  CNN_main_simple_core_core_fsm_inst_FOR_I_1_C_1_tr0 <= NOT (z_out(2));
  CNN_main_simple_core_core_fsm_inst_FOR_J_1_C_1_tr0 <= NOT (z_out(2));
  CNN_main_simple_core_core_fsm_inst_FOR_K_1_C_0_tr0 <= z_out_13(6);
  CNN_main_simple_core_core_fsm_inst_INIT_I_1_C_1_tr0 <= NOT reg_INIT_I_slc_INIT_I_acc_2_cse;
  CNN_main_simple_core_core_fsm_inst_INIT_J_1_C_0_tr0 <= NOT (z_out(2));
  CNN_main_simple_core_core_fsm_inst_INIT_L_1_C_0_tr0 <= z_out_16(5);
  CNN_main_simple_core_core_fsm_inst_FOR_B_2_C_1_tr0 <= NOT((CR1_simple_b_1_0_sva_1(0))
      XOR (CR1_simple_b_1_0_sva_1(1)));
  CNN_main_simple_core_core_fsm_inst_FOR_A_2_C_0_tr0 <= NOT((z_out_2(0)) XOR (z_out_2(1)));
  CNN_main_simple_core_core_fsm_inst_FOR_I_2_C_2_tr0 <= NOT FOR_I_2_slc_FOR_I_2_acc_2_itm;
  CNN_main_simple_core_core_fsm_inst_FOR_J_2_C_0_tr0 <= NOT (z_out(2));
  CNN_main_simple_core_core_fsm_inst_FOR_K_2_C_0_tr0 <= z_out_13(6);
  CNN_main_simple_core_core_fsm_inst_BIAS_I_1_C_2_tr0 <= NOT BIAS_I_1_slc_BIAS_I_1_acc_2_itm;
  CNN_main_simple_core_core_fsm_inst_BIAS_J_1_C_0_tr0 <= NOT (z_out(2));
  CNN_main_simple_core_core_fsm_inst_FOR_L_1_C_0_tr0 <= z_out_16(5);
  CNN_main_simple_core_core_fsm_inst_FOR_A_3_C_1_tr0 <= NOT((CR1_simple_b_1_0_sva_1(0))
      XOR (CR1_simple_b_1_0_sva_1(1)));
  CNN_main_simple_core_core_fsm_inst_FOR_B_3_C_1_tr0 <= NOT((CR1_simple_b_1_0_sva_1(0))
      XOR (CR1_simple_b_1_0_sva_1(1)));
  CNN_main_simple_core_core_fsm_inst_FOR_I_3_C_1_tr0 <= NOT (z_out(2));
  CNN_main_simple_core_core_fsm_inst_FOR_J_3_C_1_tr0 <= NOT (z_out(2));
  CNN_main_simple_core_core_fsm_inst_FOR_K_3_C_0_tr0 <= z_out_16(5);
  CNN_main_simple_core_core_fsm_inst_INIT_I_2_C_1_tr0 <= NOT reg_INIT_I_slc_INIT_I_acc_2_cse;
  CNN_main_simple_core_core_fsm_inst_INIT_J_2_C_0_tr0 <= NOT (z_out(2));
  CNN_main_simple_core_core_fsm_inst_INIT_L_2_C_0_tr0 <= NOT (z_out_7(3));
  CNN_main_simple_core_core_fsm_inst_FOR_B_4_C_1_tr0 <= NOT((CR1_simple_b_1_0_sva_1(0))
      XOR (CR1_simple_b_1_0_sva_1(1)));
  CNN_main_simple_core_core_fsm_inst_FOR_A_4_C_0_tr0 <= NOT((z_out_2(0)) XOR (z_out_2(1)));
  CNN_main_simple_core_core_fsm_inst_FOR_I_4_C_2_tr0 <= NOT FOR_I_4_slc_FOR_I_4_acc_2_itm;
  CNN_main_simple_core_core_fsm_inst_FOR_J_4_C_0_tr0 <= NOT (z_out(2));
  CNN_main_simple_core_core_fsm_inst_FOR_K_4_C_0_tr0 <= z_out_16(5);
  CNN_main_simple_core_core_fsm_inst_BIAS_I_2_C_2_tr0 <= NOT BIAS_I_2_slc_BIAS_I_2_acc_2_itm;
  CNN_main_simple_core_core_fsm_inst_BIAS_J_2_C_0_tr0 <= NOT (z_out(2));
  CNN_main_simple_core_core_fsm_inst_FOR_L_2_C_0_tr0 <= NOT (z_out_7(3));
  CNN_main_simple_core_core_fsm_inst_FOR_A_5_C_1_tr0 <= MP3_simple_a_1_0_sva(1);
  CNN_main_simple_core_core_fsm_inst_FOR_B_5_C_1_tr0 <= NOT((CR1_simple_b_1_0_sva_1(0))
      XOR (CR1_simple_b_1_0_sva_1(1)));
  CNN_main_simple_core_core_fsm_inst_FOR_I_5_C_1_tr0 <= NOT((z_out_2(0)) XOR (z_out_2(1)));
  CNN_main_simple_core_core_fsm_inst_FOR_J_5_C_1_tr0 <= NOT((z_out_2(0)) XOR (z_out_2(1)));
  CNN_main_simple_core_core_fsm_inst_FOR_K_5_C_0_tr0 <= NOT (z_out_7(3));
  CNN_main_simple_core_core_fsm_inst_FOR_K_6_C_2_tr0 <= NOT FOR_K_6_slc_FOR_K_6_acc_3_itm;
  CNN_main_simple_core_core_fsm_inst_FOR_J_6_C_0_tr0 <= NOT((z_out_2(0)) XOR (z_out_2(1)));
  CNN_main_simple_core_core_fsm_inst_FOR_K_7_C_1_tr0 <= NOT FOR_K_7_slc_FOR_K_7_acc_6_itm;
  CNN_main_simple_core_core_fsm_inst_FOR_J_7_C_1_tr0 <= NOT (z_out_7(3));
  CNN_main_simple_core_core_fsm_inst_for_C_0_tr0 <= NOT (z_out_7(3));

  memory_1_or_seb <= (fsm_output(68)) OR (fsm_output(63)) OR (fsm_output(42)) OR
      (fsm_output(37)) OR (fsm_output(16)) OR (fsm_output(11)) OR (fsm_output(82));
  memory_1_or_1_seb <= (fsm_output(68)) OR (fsm_output(55)) OR (fsm_output(29)) OR
      (fsm_output(3)) OR (fsm_output(63)) OR (fsm_output(42)) OR (fsm_output(37))
      OR (fsm_output(16)) OR (fsm_output(11)) OR (fsm_output(82)) OR (fsm_output(0));
  nand_cse_1 <= NOT(z_out_1_2 AND (z_out(2)));
  memory_1_nor_1_seb <= NOT((NOT((fsm_output(62)) OR (fsm_output(36)) OR (fsm_output(10))
      OR (fsm_output(67)) OR (fsm_output(41)) OR (fsm_output(15)) OR (fsm_output(74))
      OR (fsm_output(48)) OR (fsm_output(22)) OR (fsm_output(87)))) OR (nand_cse_1
      AND (fsm_output(22))) OR (nand_cse_1 AND (fsm_output(74))) OR (nand_cse_1 AND
      (fsm_output(48))));
  or_125_cse <= FOR_B_oelse_acc_tmp_13 OR FOR_B_oelse_2_acc_itm_13;
  reg_CR1_simple_l_1_6_0_sva_5_CR1_simple_l_or_cse <= (fsm_output(2)) OR (fsm_output(6));
  reg_CR1_simple_CR1_simple_aux_or_1_cse <= or_332_cse OR CONV_SL_1_1(fsm_output(9
      DOWNTO 8)/=STD_LOGIC_VECTOR'("00"));
  or_332_cse <= (fsm_output(13)) OR (fsm_output(19)) OR (fsm_output(14)) OR (fsm_output(6))
      OR (fsm_output(12));
  reg_CR2_simple_CR2_simple_aux_or_1_cse <= or_400_cse OR CONV_SL_1_1(fsm_output(35
      DOWNTO 34)/=STD_LOGIC_VECTOR'("00"));
  or_400_cse <= (fsm_output(39)) OR (fsm_output(45)) OR (fsm_output(40)) OR (fsm_output(32))
      OR (fsm_output(38));
  FOR_B_2_if_FOR_B_2_if_or_cse <= FOR_B_2_oelse_2_acc_itm_14 OR FOR_B_2_oelse_acc_tmp_14;
  reg_CR3_simple_CR3_simple_aux_or_1_cse <= or_468_cse OR CONV_SL_1_1(fsm_output(61
      DOWNTO 60)/=STD_LOGIC_VECTOR'("00"));
  or_468_cse <= (fsm_output(65)) OR (fsm_output(71)) OR (fsm_output(66)) OR (fsm_output(58))
      OR (fsm_output(64));
  FOR_B_4_if_FOR_B_4_if_or_cse <= (z_out_22(15)) OR FOR_B_4_oelse_acc_tmp_15;
  reg_MP3_simple_b_1_MP3_simple_b_or_cse <= (fsm_output(73)) OR (fsm_output(77));
  FOR_J_7_or_29_rgt <= (fsm_output(87)) OR ((NOT FOR_J_7_and_21_cse_sva) AND (fsm_output(88)));
  FOR_J_7_and_81_rgt <= FOR_J_7_and_21_cse_sva AND (fsm_output(88));
  FOR_J_7_or_2_rgt <= (fsm_output(87)) OR ((NOT FOR_J_7_and_20_cse_sva) AND (fsm_output(88)));
  FOR_J_7_and_27_rgt <= FOR_J_7_and_20_cse_sva AND (fsm_output(88));
  FOR_J_7_or_26_rgt <= (fsm_output(87)) OR ((NOT FOR_J_7_and_19_cse_sva) AND (fsm_output(88)));
  FOR_J_7_and_75_rgt <= FOR_J_7_and_19_cse_sva AND (fsm_output(88));
  FOR_J_7_or_23_rgt <= (fsm_output(87)) OR ((NOT FOR_J_7_and_18_cse_sva) AND (fsm_output(88)));
  FOR_J_7_and_69_rgt <= FOR_J_7_and_18_cse_sva AND (fsm_output(88));
  FOR_J_7_or_20_rgt <= (fsm_output(87)) OR ((NOT FOR_J_7_and_17_cse_sva) AND (fsm_output(88)));
  FOR_J_7_and_63_rgt <= FOR_J_7_and_17_cse_sva AND (fsm_output(88));
  FOR_J_7_or_17_rgt <= (fsm_output(87)) OR ((NOT FOR_J_7_and_16_cse_sva) AND (fsm_output(88)));
  FOR_J_7_and_57_rgt <= FOR_J_7_and_16_cse_sva AND (fsm_output(88));
  FOR_J_7_or_14_rgt <= (fsm_output(87)) OR ((NOT FOR_J_7_and_15_cse_sva) AND (fsm_output(88)));
  FOR_J_7_and_51_rgt <= FOR_J_7_and_15_cse_sva AND (fsm_output(88));
  FOR_J_7_or_11_rgt <= (fsm_output(87)) OR ((NOT FOR_J_7_and_14_cse_sva) AND (fsm_output(88)));
  FOR_J_7_and_45_rgt <= FOR_J_7_and_14_cse_sva AND (fsm_output(88));
  FOR_J_7_or_8_rgt <= (fsm_output(87)) OR ((NOT FOR_J_7_and_13_cse_sva) AND (fsm_output(88)));
  FOR_J_7_and_39_rgt <= FOR_J_7_and_13_cse_sva AND (fsm_output(88));
  FOR_J_7_or_5_rgt <= (fsm_output(87)) OR ((NOT FOR_J_7_and_12_cse_sva) AND (fsm_output(88)));
  FOR_J_7_and_33_rgt <= FOR_J_7_and_12_cse_sva AND (fsm_output(88));
  CR1_simple_aux_15_lpi_7_mx1 <= MUX_s_1_2_2((FOR_B_if_acc_psp_sva_1(18)), CR1_simple_aux_15_lpi_7,
      FOR_B_lor_2_lpi_7_dfm_st);
  FOR_B_if_nor_2_nl <= NOT(MUX_v_14_2_2((FOR_B_if_acc_psp_sva_1(14 DOWNTO 1)), STD_LOGIC_VECTOR'("11111111111111"),
      FOR_B_if_nor_ovfl_sva_1));
  FOR_B_if_FOR_B_if_nor_nl <= NOT(MUX_v_14_2_2(FOR_B_if_nor_2_nl, STD_LOGIC_VECTOR'("11111111111111"),
      FOR_B_if_and_unfl_sva_1));
  CR1_simple_aux_14_1_lpi_7_mx1 <= MUX_v_14_2_2(FOR_B_if_FOR_B_if_nor_nl, CR1_simple_aux_14_1_lpi_7,
      FOR_B_lor_2_lpi_7_dfm_st);
  FOR_B_if_FOR_B_if_nor_1_nl <= NOT((NOT((FOR_B_if_acc_psp_sva_1(0)) OR FOR_B_if_nor_ovfl_sva_1))
      OR FOR_B_if_and_unfl_sva_1);
  CR1_simple_aux_0_lpi_7_mx1 <= MUX_s_1_2_2(FOR_B_if_FOR_B_if_nor_1_nl, CR1_simple_aux_0_lpi_7,
      FOR_B_lor_2_lpi_7_dfm_st);
  FOR_B_if_acc_10_psp_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_SIGNED(SIGNED(FOR_B_if_acc_5_sdt_1(5
      DOWNTO 1)), 5), 7) + CONV_UNSIGNED(CONV_SIGNED(SIGNED(FOR_B_acc_1_psp_sva_1),
      6), 7), 7));
  FOR_B_if_acc_5_sdt_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(FOR_B_acc_1_psp_sva_1)
      + CONV_SIGNED(CONV_SIGNED(SIGNED(z_out_16(5 DOWNTO 3)), 3), 6), 6));
  FOR_B_acc_1_psp_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_SIGNED(SIGNED(z_out_15_1_0),
      2), 6) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(CR1_simple_i_2_4_0_sva), 5), 6),
      6));
  FOR_B_oelse_2_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(NOT
      (z_out_16(5 DOWNTO 3))),13))) + UNSIGNED'( "00000000000011"), 14));
  FOR_B_oelse_2_acc_itm_13 <= READSLICE_1_14(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(FOR_B_oelse_2_acc_nl),
      14)), 13);
  FOR_B_oelse_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(NOT
      (FOR_B_acc_1_psp_sva_1(5 DOWNTO 3))),13))) + UNSIGNED'( "00000000000011"),
      14));
  FOR_B_oelse_acc_tmp_13 <= READSLICE_1_14(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(FOR_B_oelse_acc_nl),
      14)), 13);
  FOR_B_if_acc_psp_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_SIGNED(SIGNED(CR1_simple_aux_15_lpi_7
      & CR1_simple_aux_14_1_lpi_7 & CR1_simple_aux_0_lpi_7), 16), 19) + UNSIGNED(z_out_18_31_12(19
      DOWNTO 1)), 19));
  FOR_B_if_nor_ovfl_sva_1 <= NOT((FOR_B_if_acc_psp_sva_1(18)) OR (NOT(CONV_SL_1_1(FOR_B_if_acc_psp_sva_1(17
      DOWNTO 15)/=STD_LOGIC_VECTOR'("000")))));
  FOR_B_if_and_unfl_sva_1 <= (FOR_B_if_acc_psp_sva_1(18)) AND (NOT(CONV_SL_1_1(FOR_B_if_acc_psp_sva_1(17
      DOWNTO 15)=STD_LOGIC_VECTOR'("111"))));
  FOR_I_nor_2_cse <= NOT(CONV_SL_1_1(z_out_22(16 DOWNTO 15)/=STD_LOGIC_VECTOR'("01")));
  FOR_I_and_4_cse <= CONV_SL_1_1(z_out_22(16 DOWNTO 15)=STD_LOGIC_VECTOR'("10"));
  or_141_cse <= reg_FOR_A_1_lor_lpi_6_dfm_cse OR (NOT (z_out_22(16)));
  MP1_simple_bigger_lpi_6_mx1 <= MUX_v_16_2_2(memory_1_rsci_q_d, MP1_simple_bigger_lpi_6,
      or_141_cse);
  FOR_A_1_oelse_acc_1_ncse_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MP1_simple_i_4_1_sva)
      + CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(MP1_simple_a_1_0_sva(1), 1), 1),
      4), 4));
  FOR_B_1_if_acc_3_sdt_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(MP1_simple_k_6_0_sva_5_0),
      6), 7) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(z_out_23(4 DOWNTO 1)), 4), 7),
      7));
  CR2_simple_aux_15_lpi_7_mx1 <= MUX_s_1_2_2((z_out_24(19)), CR2_simple_aux_15_lpi_7,
      FOR_B_2_lor_2_lpi_7_dfm_st);
  FOR_B_2_if_nor_2_nl <= NOT(MUX_v_14_2_2((z_out_24(14 DOWNTO 1)), STD_LOGIC_VECTOR'("11111111111111"),
      FOR_B_2_if_nor_ovfl_sva_1));
  FOR_B_2_if_FOR_B_2_if_nor_cse <= NOT(MUX_v_14_2_2(FOR_B_2_if_nor_2_nl, STD_LOGIC_VECTOR'("11111111111111"),
      FOR_B_2_if_and_unfl_sva_1));
  CR2_simple_aux_14_1_lpi_7_mx1 <= MUX_v_14_2_2(FOR_B_2_if_FOR_B_2_if_nor_cse, CR2_simple_aux_14_1_lpi_7,
      FOR_B_2_lor_2_lpi_7_dfm_st);
  FOR_B_2_if_FOR_B_2_if_nor_1_cse <= NOT((NOT((z_out_24(0)) OR FOR_B_2_if_nor_ovfl_sva_1))
      OR FOR_B_2_if_and_unfl_sva_1);
  CR2_simple_aux_0_lpi_7_mx1 <= MUX_s_1_2_2(FOR_B_2_if_FOR_B_2_if_nor_1_cse, CR2_simple_aux_0_lpi_7,
      FOR_B_2_lor_2_lpi_7_dfm_st);
  FOR_B_2_if_acc_8_sdt_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(CR2_simple_k_6_0_sva_5_0_1),
      6), 7) + CONV_UNSIGNED(CONV_SIGNED(SIGNED(FOR_B_2_if_acc_9_psp_1(5 DOWNTO 1)),
      5), 7), 7));
  FOR_B_2_if_acc_9_psp_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_SIGNED(SIGNED(z_out_16(4
      DOWNTO 1)), 4), 6) + CONV_UNSIGNED(CONV_SIGNED(SIGNED(FOR_B_2_acc_1_psp_sva_1),
      5), 6), 6));
  CR2_simple_j_aux_4_0_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_SIGNED(SIGNED(z_out_14_1_0),
      2), 5) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(CR2_simple_j_2_3_0_sva), 4),
      5), 5));
  FOR_B_2_acc_1_psp_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_SIGNED(SIGNED(z_out_15_1_0),
      2), 5) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(CR2_simple_i_2_3_0_sva), 4), 5),
      5));
  FOR_B_2_oelse_2_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(NOT
      (CR2_simple_j_aux_4_0_sva_1(4 DOWNTO 2))),14))) + UNSIGNED'( "000000000000011"),
      15));
  FOR_B_2_oelse_2_acc_itm_14 <= READSLICE_1_15(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(FOR_B_2_oelse_2_acc_nl),
      15)), 14);
  FOR_B_2_oelse_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(NOT
      (FOR_B_2_acc_1_psp_sva_1(4 DOWNTO 2))),14))) + UNSIGNED'( "000000000000011"),
      15));
  FOR_B_2_oelse_acc_tmp_14 <= READSLICE_1_15(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(FOR_B_2_oelse_acc_nl),
      15)), 14);
  FOR_B_2_if_nor_ovfl_sva_1 <= NOT((z_out_24(19)) OR (NOT(CONV_SL_1_1(z_out_24(18
      DOWNTO 15)/=STD_LOGIC_VECTOR'("0000")))));
  FOR_B_2_if_and_unfl_sva_1 <= (z_out_24(19)) AND (NOT(CONV_SL_1_1(z_out_24(18 DOWNTO
      15)=STD_LOGIC_VECTOR'("1111"))));
  MP2_simple_bigger_lpi_6_mx1 <= MUX_v_16_2_2(memory_1_rsci_q_d, MP2_simple_bigger_lpi_6,
      or_141_cse);
  FOR_A_3_oelse_acc_1_ncse_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MP2_simple_i_3_1_sva)
      + CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(MP2_simple_a_1_0_sva(1), 1), 1),
      3), 3));
  FOR_B_3_if_acc_sdt_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MP2_simple_j_N_2_0_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(MP2_simple_i_N_2_0_sva_1(2 DOWNTO 1)),
      2), 3), 3));
  INIT_I_2_acc_6_sdt_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(CR3_simple_l_1_4_0_sva)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(z_out_26), 4), 5), 5));
  CR3_simple_aux_15_lpi_7_mx1 <= MUX_s_1_2_2((z_out_24(19)), CR3_simple_aux_15_lpi_7,
      FOR_B_4_lor_2_lpi_7_dfm_st);
  CR3_simple_aux_14_1_lpi_7_mx1 <= MUX_v_14_2_2(FOR_B_2_if_FOR_B_2_if_nor_cse, CR3_simple_aux_14_1_lpi_7,
      FOR_B_4_lor_2_lpi_7_dfm_st);
  CR3_simple_aux_0_lpi_7_mx1 <= MUX_s_1_2_2(FOR_B_2_if_FOR_B_2_if_nor_1_cse, CR3_simple_aux_0_lpi_7,
      FOR_B_4_lor_2_lpi_7_dfm_st);
  FOR_B_4_if_acc_12_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_SIGNED(SIGNED(FOR_B_4_if_acc_6_sdt_1(4
      DOWNTO 1)), 4), 5) + CONV_SIGNED(CONV_SIGNED(SIGNED(FOR_B_4_acc_1_psp_1_sva_1),
      4), 5), 5));
  FOR_B_4_if_acc_11_sdt_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(SIGNED(FOR_B_4_if_acc_12_nl),
      7) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(CR3_simple_k_5_0_sva_4_0), 5), 7),
      7));
  FOR_B_4_if_acc_6_sdt_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_SIGNED(SIGNED(FOR_B_4_acc_1_psp_1_sva_1),
      4), 5) + CONV_SIGNED(CONV_SIGNED(SIGNED(CR3_simple_j_aux_3_0_sva_1(3 DOWNTO
      1)), 3), 5), 5));
  CR3_simple_j_aux_3_0_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_SIGNED(SIGNED(z_out_15_1_0),
      2), 4) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(CR3_simple_j_2_2_0_sva), 3),
      4), 4));
  FOR_B_4_acc_1_psp_1_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_SIGNED(SIGNED(z_out_14_1_0),
      2), 4) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(CR3_simple_i_2_2_0_sva), 3), 4),
      4));
  FOR_B_4_if_acc_9_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_SIGNED(SIGNED(z_out),
      3), 4) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(z_out_10(5 DOWNTO 3)), 3), 4),
      4));
  FOR_B_4_if_acc_10_sdt_4_0_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(SIGNED(FOR_B_4_if_acc_9_nl),
      5) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(CR3_simple_b_1_0_sva & STD_LOGIC_VECTOR'(
      "01")), 4), 5), 5));
  FOR_B_4_oelse_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(NOT
      (FOR_B_4_acc_1_psp_1_sva_1(3 DOWNTO 1))),15))) + UNSIGNED'( "0000000000000011"),
      16));
  FOR_B_4_oelse_acc_tmp_15 <= READSLICE_1_16(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(FOR_B_4_oelse_acc_nl),
      16)), 15);
  MP3_simple_bigger_lpi_6_mx1 <= MUX_v_16_2_2(memory_1_rsci_q_d, MP3_simple_bigger_lpi_6,
      or_141_cse);
  FOR_J_7_and_stg_2_1_sva_1 <= FOR_J_7_and_stg_1_1_sva_1 AND (NOT (perceptron_simple_j_3_0_sva(2)));
  FOR_J_7_and_stg_2_0_sva_1 <= FOR_J_7_and_stg_1_0_sva_1 AND (NOT (perceptron_simple_j_3_0_sva(2)));
  FOR_J_7_and_stg_1_3_sva_1 <= CONV_SL_1_1(perceptron_simple_j_3_0_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  FOR_J_7_and_stg_1_2_sva_1 <= CONV_SL_1_1(perceptron_simple_j_3_0_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"));
  FOR_J_7_and_stg_1_1_sva_1 <= CONV_SL_1_1(perceptron_simple_j_3_0_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"));
  FOR_J_7_and_stg_1_0_sva_1 <= NOT(CONV_SL_1_1(perceptron_simple_j_3_0_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("00")));
  perceptron_simple_k_7_0_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(perceptron_simple_k_7_0_sva)
      + UNSIGNED'( "00000001"), 8));
  FOR_K_7_acc_8_sdt_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(perceptron_simple_k_7_0_sva)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(perceptron_simple_j_3_0_sva(3 DOWNTO
      1)), 3), 8), 8));
  FOR_K_7_acc_7_psp_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_SIGNED(SIGNED(FOR_K_7_mux_28_itm
      & FOR_K_7_mux_29_itm & FOR_K_7_mux_30_itm), 16), 17) + UNSIGNED(z_out_18_31_12(19
      DOWNTO 3)), 17));
  FOR_K_7_FOR_K_7_nor_2_psp_sva_1 <= NOT((NOT((FOR_K_7_acc_7_psp_sva_1(0)) OR FOR_K_7_nor_ovfl_sva_1))
      OR FOR_K_7_and_unfl_sva_1);
  FOR_K_7_nor_3_nl <= NOT(MUX_v_14_2_2((FOR_K_7_acc_7_psp_sva_1(14 DOWNTO 1)), STD_LOGIC_VECTOR'("11111111111111"),
      FOR_K_7_nor_ovfl_sva_1));
  FOR_K_7_FOR_K_7_nor_1_psp_sva_1 <= NOT(MUX_v_14_2_2(FOR_K_7_nor_3_nl, STD_LOGIC_VECTOR'("11111111111111"),
      FOR_K_7_and_unfl_sva_1));
  FOR_K_7_nor_ovfl_sva_1 <= NOT(CONV_SL_1_1(FOR_K_7_acc_7_psp_sva_1(16 DOWNTO 15)/=STD_LOGIC_VECTOR'("01")));
  FOR_K_7_and_unfl_sva_1 <= CONV_SL_1_1(FOR_K_7_acc_7_psp_sva_1(16 DOWNTO 15)=STD_LOGIC_VECTOR'("10"));
  max_sva_14_1_mx1 <= MUX_v_14_2_2(max_sva_14_1, for_slc_Prob_16_15_0_cse_sva_14_1_1,
      z_out_22(16));
  for_slc_Prob_16_15_0_cse_sva_14_1_1 <= MUX_v_14_10_2(Prob_0_sva_2_14_1, Prob_1_14_1_sva_2,
      Prob_2_14_1_sva_2, Prob_3_14_1_sva_2, Prob_4_14_1_sva_2, Prob_5_14_1_sva_2,
      Prob_6_14_1_sva_2, Prob_7_14_1_sva_2, Prob_8_14_1_sva_2, Prob_9_14_1_sva_2,
      k_sva);
  for_slc_Prob_16_15_0_cse_sva_15_1 <= MUX_s_1_10_2(Prob_0_sva_2_15, Prob_1_15_sva_2,
      Prob_2_15_sva_2, Prob_3_15_sva_2, Prob_4_15_sva_2, Prob_5_15_sva_2, Prob_6_15_sva_2,
      Prob_7_15_sva_2, Prob_8_15_sva_2, Prob_9_15_sva_2, k_sva);
  for_slc_Prob_16_15_0_cse_sva_0_1 <= MUX_s_1_10_2(Prob_0_sva_2_0, Prob_1_0_sva_2,
      Prob_2_0_sva_2, Prob_3_0_sva_2, Prob_4_0_sva_2, Prob_5_0_sva_2, Prob_6_0_sva_2,
      Prob_7_0_sva_2, Prob_8_0_sva_2, Prob_9_0_sva_2, k_sva);
  FOR_I_6_FOR_I_6_xnor_cse <= NOT((z_out_2(0)) XOR (z_out_2(1)));
  and_4_cse <= CONV_SL_1_1(fsm_output(10 DOWNTO 9)/=STD_LOGIC_VECTOR'("00"));
  and_10_cse <= CONV_SL_1_1(fsm_output(36 DOWNTO 35)/=STD_LOGIC_VECTOR'("00"));
  and_16_cse <= CONV_SL_1_1(fsm_output(62 DOWNTO 61)/=STD_LOGIC_VECTOR'("00"));
  or_dcpl_53 <= (fsm_output(1)) OR (fsm_output(91));
  and_dcpl_6 <= NOT((fsm_output(76)) OR (fsm_output(50)));
  and_dcpl_133 <= CONV_SL_1_1(perceptron_simple_j_3_0_sva(3 DOWNTO 2)=STD_LOGIC_VECTOR'("10"));
  or_dcpl_130 <= CONV_SL_1_1(perceptron_simple_j_3_0_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"));
  or_dcpl_131 <= CONV_SL_1_1(perceptron_simple_j_3_0_sva(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("10"));
  and_dcpl_136 <= NOT(CONV_SL_1_1(perceptron_simple_j_3_0_sva(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")));
  or_dcpl_134 <= CONV_SL_1_1(perceptron_simple_j_3_0_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"));
  or_dcpl_135 <= CONV_SL_1_1(perceptron_simple_j_3_0_sva(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"));
  and_dcpl_141 <= CONV_SL_1_1(perceptron_simple_j_3_0_sva(3 DOWNTO 2)=STD_LOGIC_VECTOR'("01"));
  or_dcpl_139 <= NOT(CONV_SL_1_1(perceptron_simple_j_3_0_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")));
  or_dcpl_140 <= CONV_SL_1_1(perceptron_simple_j_3_0_sva(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"));
  or_dcpl_142 <= CONV_SL_1_1(perceptron_simple_j_3_0_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"));
  and_285_cse <= (NOT(FOR_B_2_oelse_acc_tmp_14 OR FOR_B_2_oelse_2_acc_itm_14)) AND
      (fsm_output(33));
  and_283_cse <= (NOT(FOR_B_4_oelse_acc_tmp_15 OR (z_out_22(15)))) AND (fsm_output(59));
  and_307_cse <= FOR_B_2_if_FOR_B_2_if_or_cse AND (fsm_output(33));
  and_316_cse <= z_out_1_2 AND (z_out(2)) AND (fsm_output(22));
  and_318_cse <= z_out_1_2 AND (z_out(2)) AND (fsm_output(48));
  and_317_cse <= z_out_1_2 AND (z_out(2)) AND (fsm_output(74));
  and_386_cse <= (z_out_7(3)) AND (fsm_output(89));
  or_tmp_111 <= (NOT((fsm_output(33)) OR (fsm_output(0)))) OR and_307_cse;
  or_tmp_117 <= (NOT(FOR_B_oelse_acc_tmp_13 OR FOR_B_oelse_2_acc_itm_13)) AND (fsm_output(7));
  or_tmp_125 <= NOT(CONV_SL_1_1(fsm_output(88 DOWNTO 86)/=STD_LOGIC_VECTOR'("000")));
  or_tmp_376 <= CONV_SL_1_1(fsm_output(90 DOWNTO 89)/=STD_LOGIC_VECTOR'("00"));
  or_tmp_379 <= and_dcpl_133 AND FOR_J_7_and_stg_1_1_sva_1 AND (fsm_output(86));
  or_tmp_380 <= (or_dcpl_131 OR or_dcpl_130) AND (fsm_output(86));
  or_tmp_383 <= CONV_SL_1_1(fsm_output(88 DOWNTO 87)/=STD_LOGIC_VECTOR'("00"));
  or_tmp_392 <= and_dcpl_136 AND FOR_J_7_and_stg_1_0_sva_1 AND (fsm_output(86));
  or_tmp_393 <= (or_dcpl_135 OR or_dcpl_134) AND (fsm_output(86));
  or_tmp_405 <= and_dcpl_133 AND FOR_J_7_and_stg_1_0_sva_1 AND (fsm_output(86));
  or_tmp_406 <= (or_dcpl_131 OR or_dcpl_134) AND (fsm_output(86));
  or_tmp_418 <= and_dcpl_136 AND FOR_J_7_and_stg_1_1_sva_1 AND (fsm_output(86));
  or_tmp_419 <= (or_dcpl_135 OR or_dcpl_130) AND (fsm_output(86));
  or_tmp_431 <= and_dcpl_141 AND FOR_J_7_and_stg_1_3_sva_1 AND (fsm_output(86));
  or_tmp_432 <= (or_dcpl_140 OR or_dcpl_139) AND (fsm_output(86));
  or_tmp_444 <= and_dcpl_136 AND FOR_J_7_and_stg_1_2_sva_1 AND (fsm_output(86));
  or_tmp_445 <= (or_dcpl_135 OR or_dcpl_142) AND (fsm_output(86));
  or_tmp_457 <= and_dcpl_141 AND FOR_J_7_and_stg_1_2_sva_1 AND (fsm_output(86));
  or_tmp_458 <= (or_dcpl_140 OR or_dcpl_142) AND (fsm_output(86));
  or_tmp_470 <= and_dcpl_136 AND FOR_J_7_and_stg_1_3_sva_1 AND (fsm_output(86));
  or_tmp_471 <= (or_dcpl_135 OR or_dcpl_139) AND (fsm_output(86));
  or_tmp_483 <= and_dcpl_141 AND FOR_J_7_and_stg_1_1_sva_1 AND (fsm_output(86));
  or_tmp_484 <= (or_dcpl_140 OR or_dcpl_130) AND (fsm_output(86));
  or_tmp_496 <= and_dcpl_141 AND FOR_J_7_and_stg_1_0_sva_1 AND (fsm_output(86));
  or_tmp_497 <= (or_dcpl_140 OR or_dcpl_134) AND (fsm_output(86));
  memory_2_rsci_wadr_d_mx0c0 <= and_dcpl_6 AND (NOT (fsm_output(24)));
  memory_2_rsci_radr_d_mx0c0 <= (NOT((fsm_output(81)) OR (fsm_output(59)) OR (fsm_output(33))))
      OR (FOR_B_4_if_FOR_B_4_if_or_cse AND (fsm_output(59))) OR and_307_cse;
  reshape_simple_add_N_10_0_lpi_4_mx0c1 <= CONV_SL_1_1(fsm_output(85 DOWNTO 83)/=STD_LOGIC_VECTOR'("000"));
  INIT_I_asn_CR1_simple_add_AF_10_INIT_I_acc_sdt <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(z_out_17
      & (z_out_10(4 DOWNTO 2))) + UNSIGNED(CR1_simple_l_1_6_0_sva_5_0(4 DOWNTO 0)),
      5));
  or_220_ssc <= (fsm_output(82)) OR (fsm_output(0));
  FOR_A_1_if_asn_MP1_simple_add_M_10_FOR_A_1_if_acc_sdt <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(z_out_17
      & (z_out_23(3 DOWNTO 1))) + UNSIGNED(MP1_simple_k_6_0_sva_5_0(4 DOWNTO 0)),
      5));
  FOR_B_if_asn_CR1_simple_add_M_10_FOR_B_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(CR1_simple_k_1_0_sva
      & '0' & CR1_simple_k_1_0_sva) + UNSIGNED(FOR_B_if_acc_10_psp_1(6 DOWNTO 2)),
      5));
  BIAS_I_BIAS_I_and_2_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(FOR_B_if_asn_CR1_simple_add_M_10_FOR_B_if_acc_nl),
      5)), or_tmp_117);
  FOR_K_FOR_K_and_5_nl <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), (FOR_B_if_acc_10_psp_1(1
      DOWNTO 0)), or_tmp_117);
  BIAS_I_BIAS_I_and_3_nl <= (FOR_B_if_acc_5_sdt_1(0)) AND or_tmp_117;
  BIAS_I_2_BIAS_I_2_and_3_nl <= MUX_v_3_2_2(STD_LOGIC_VECTOR'("000"), (z_out_16(2
      DOWNTO 0)), or_tmp_117);
  image_rsci_radr_d <= BIAS_I_BIAS_I_and_2_nl & FOR_K_FOR_K_and_5_nl & BIAS_I_BIAS_I_and_3_nl
      & BIAS_I_2_BIAS_I_2_and_3_nl;
  image_rsci_re_d_pff <= or_tmp_117;
  FOR_K_FOR_K_and_4_nl <= (((z_out_7(3)) AND (CR1_simple_a_1_0_sva(0))) XOR (CR1_simple_a_1_0_sva(1)))
      AND or_tmp_117;
  FOR_K_FOR_K_and_11_nl <= ((z_out_7(3)) XOR (CR1_simple_a_1_0_sva(0))) AND or_tmp_117;
  BIAS_I_2_BIAS_I_2_and_2_nl <= MUX_v_3_2_2(STD_LOGIC_VECTOR'("000"), (z_out_7(2
      DOWNTO 0)), or_tmp_117);
  CR1_simple_l_nor_nl <= NOT((NOT((fsm_output(7)) OR (fsm_output(0)))) OR (or_125_cse
      AND (fsm_output(7))));
  CR1_simple_l_CR1_simple_l_and_1_nl <= MUX_v_6_2_2(STD_LOGIC_VECTOR'("000000"),
      CR1_simple_l_6_0_sva_5_0_1, CR1_simple_l_nor_nl);
  F_1_rsci_radr_d <= FOR_K_FOR_K_and_4_nl & FOR_K_FOR_K_and_11_nl & BIAS_I_2_BIAS_I_2_and_2_nl
      & CR1_simple_l_CR1_simple_l_and_1_nl;
  B_1_nor_nl <= NOT((NOT((fsm_output(17)) OR (fsm_output(18)) OR (fsm_output(14))
      OR (fsm_output(0)))) OR ((NOT BIAS_I_slc_BIAS_I_acc_2_itm) AND (fsm_output(17)))
      OR (((z_out_2(0)) XOR (z_out_2(1))) AND (fsm_output(14))) OR ((NOT (z_out(2)))
      AND (fsm_output(18))));
  B_1_rsci_radr_d <= MUX_v_6_2_2(STD_LOGIC_VECTOR'("000000"), CR1_simple_l_6_0_sva_5_0_1,
      B_1_nor_nl);
  B_1_rsci_re_d <= (BIAS_I_slc_BIAS_I_acc_2_itm AND (fsm_output(17))) OR (FOR_I_6_FOR_I_6_xnor_cse
      AND (fsm_output(14))) OR ((z_out(2)) AND (fsm_output(18)));
  BIAS_I_2_BIAS_I_2_and_1_nl <= MUX_v_3_2_2(STD_LOGIC_VECTOR'("000"), z_out_3, and_285_cse);
  BIAS_I_BIAS_I_and_1_nl <= (z_out_4(0)) AND and_285_cse;
  CR2_simple_k_not_nl <= NOT or_tmp_111;
  CR2_simple_k_CR2_simple_k_and_nl <= MUX_v_6_2_2(STD_LOGIC_VECTOR'("000000"), CR2_simple_k_6_0_sva_5_0_1,
      CR2_simple_k_not_nl);
  CR2_simple_l_not_nl <= NOT or_tmp_111;
  CR2_simple_l_CR2_simple_l_and_1_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), CR2_simple_l_5_0_sva_4_0_1,
      CR2_simple_l_not_nl);
  F_2_rsci_radr_d <= BIAS_I_2_BIAS_I_2_and_1_nl & BIAS_I_BIAS_I_and_1_nl & CR2_simple_k_CR2_simple_k_and_nl
      & CR2_simple_l_CR2_simple_l_and_1_nl;
  F_2_rsci_re_d <= and_285_cse;
  B_2_nor_nl <= NOT((NOT((fsm_output(43)) OR (fsm_output(44)) OR (fsm_output(40))
      OR (fsm_output(0)))) OR ((NOT BIAS_I_1_slc_BIAS_I_1_acc_2_itm) AND (fsm_output(43)))
      OR ((NOT (z_out(2))) AND (fsm_output(44))) OR ((NOT (z_out_13(6))) AND (fsm_output(40))));
  B_2_rsci_radr_d <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), CR2_simple_l_5_0_sva_4_0_1,
      B_2_nor_nl);
  B_2_rsci_re_d <= (BIAS_I_1_slc_BIAS_I_1_acc_2_itm AND (fsm_output(43))) OR ((z_out(2))
      AND (fsm_output(44))) OR ((z_out_13(6)) AND (fsm_output(40)));
  FOR_K_FOR_K_and_3_nl <= (((FOR_B_4_if_acc_10_sdt_4_0_1(4)) AND (CR3_simple_a_1_0_sva(0)))
      XOR (FOR_B_4_if_acc_10_sdt_4_0_1(4)) XOR (CR3_simple_a_1_0_sva(1))) AND and_283_cse;
  FOR_K_FOR_K_and_10_nl <= ((FOR_B_4_if_acc_10_sdt_4_0_1(4)) XOR (CR3_simple_a_1_0_sva(0)))
      AND and_283_cse;
  BIAS_I_1_BIAS_I_1_and_nl <= MUX_v_4_2_2(STD_LOGIC_VECTOR'("0000"), (FOR_B_4_if_acc_10_sdt_4_0_1(3
      DOWNTO 0)), and_283_cse);
  BIAS_I_2_BIAS_I_2_and_nl <= MUX_v_3_2_2(STD_LOGIC_VECTOR'("000"), (z_out_10(2 DOWNTO
      0)), and_283_cse);
  FOR_K_FOR_K_and_2_nl <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), (z_out_11(1 DOWNTO
      0)), and_283_cse);
  FOR_K_FOR_K_and_1_nl <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), (CR3_simple_l_4_0_sva(1
      DOWNTO 0)), and_283_cse);
  F_3_rsci_radr_d <= FOR_K_FOR_K_and_3_nl & FOR_K_FOR_K_and_10_nl & BIAS_I_1_BIAS_I_1_and_nl
      & BIAS_I_2_BIAS_I_2_and_nl & FOR_K_FOR_K_and_2_nl & FOR_K_FOR_K_and_1_nl;
  F_3_rsci_re_d <= and_283_cse;
  B_3_nor_nl <= NOT((NOT((fsm_output(69)) OR (fsm_output(70)) OR (fsm_output(66))
      OR (fsm_output(0)))) OR ((NOT BIAS_I_2_slc_BIAS_I_2_acc_2_itm) AND (fsm_output(69)))
      OR ((NOT (z_out(2))) AND (fsm_output(70))) OR ((NOT (z_out_16(5))) AND (fsm_output(66))));
  B_3_rsci_radr_d <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), CR3_simple_l_4_0_sva,
      B_3_nor_nl);
  B_3_rsci_re_d <= (BIAS_I_2_slc_BIAS_I_2_acc_2_itm AND (fsm_output(69))) OR ((z_out(2))
      AND (fsm_output(70))) OR ((z_out_16(5)) AND (fsm_output(66)));
  FOR_K_7_acc_9_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(FOR_K_7_acc_8_sdt_1(7
      DOWNTO 2)), 6), 8) + UNSIGNED(perceptron_simple_k_7_0_sva), 8));
  FOR_K_7_FOR_K_7_and_nl <= MUX_v_8_2_2(STD_LOGIC_VECTOR'("00000000"), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(FOR_K_7_acc_9_nl),
      8)), (fsm_output(87)));
  FOR_K_FOR_K_and_nl <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), (FOR_K_7_acc_8_sdt_1(1
      DOWNTO 0)), (fsm_output(87)));
  BIAS_I_BIAS_I_and_nl <= (perceptron_simple_j_3_0_sva(0)) AND (fsm_output(87));
  P_W_rsci_radr_d <= FOR_K_7_FOR_K_7_and_nl & FOR_K_FOR_K_and_nl & BIAS_I_BIAS_I_and_nl;
  P_W_rsci_re_d <= fsm_output(87);
  P_B_rsci_radr_d <= MUX_v_4_2_2(STD_LOGIC_VECTOR'("0000"), z_out_5, and_386_cse);
  P_B_rsci_re_d <= (FOR_I_6_FOR_I_6_xnor_cse AND (fsm_output(85))) OR and_386_cse;
  memory_1_or_2_cse <= (fsm_output(10)) OR (fsm_output(15));
  memory_1_or_5_cse <= (fsm_output(36)) OR (fsm_output(41));
  memory_1_or_6_cse_1 <= (fsm_output(62)) OR (fsm_output(67));
  memory_1_or_3_cse <= (fsm_output(36)) OR (fsm_output(41)) OR and_318_cse;
  memory_1_or_12_cse <= (fsm_output(62)) OR (fsm_output(67)) OR and_317_cse;
  memory_1_or_13_cse <= (fsm_output(10)) OR (fsm_output(15)) OR (fsm_output(36))
      OR (fsm_output(41)) OR and_318_cse;
  memory_1_mux1h_1_nl <= MUX1HOT_s_1_3_2((z_out_19(4)), (FOR_A_1_if_asn_MP1_simple_add_M_10_FOR_A_1_if_acc_sdt(4)),
      (z_out_7(3)), STD_LOGIC_VECTOR'( memory_1_or_2_cse & and_316_cse & memory_1_or_3_cse));
  memory_1_and_1_nl <= memory_1_mux1h_1_nl AND (NOT((fsm_output(62)) OR (fsm_output(67))
      OR and_317_cse OR (fsm_output(87)))) AND memory_1_nor_1_seb;
  memory_1_mux1h_5_nl <= MUX1HOT_v_4_5_2((z_out_19(3 DOWNTO 0)), (FOR_A_1_if_asn_MP1_simple_add_M_10_FOR_A_1_if_acc_sdt(3
      DOWNTO 0)), ((z_out_7(2 DOWNTO 0)) & (z_out_10(2))), (z_out_12(4 DOWNTO 1)),
      (STD_LOGIC_VECTOR'( "00") & (perceptron_simple_k_7_0_sva(7 DOWNTO 6))), STD_LOGIC_VECTOR'(
      memory_1_or_2_cse & and_316_cse & memory_1_or_3_cse & memory_1_or_12_cse &
      (fsm_output(87))));
  memory_1_mux1h_12_nl <= MUX1HOT_s_1_4_2((z_out_10(1)), (z_out_23(0)), (z_out_12(0)),
      (perceptron_simple_k_7_0_sva(5)), STD_LOGIC_VECTOR'( memory_1_or_13_cse & and_316_cse
      & memory_1_or_12_cse & (fsm_output(87))));
  memory_1_mux1h_13_nl <= MUX1HOT_s_1_5_2((z_out_10(0)), (z_out_8(0)), (z_out_20(2)),
      (z_out_21(2)), (perceptron_simple_k_7_0_sva(4)), STD_LOGIC_VECTOR'( memory_1_or_13_cse
      & and_316_cse & memory_1_or_6_cse_1 & and_317_cse & (fsm_output(87))));
  memory_1_and_4_nl <= MUX_v_6_2_2(STD_LOGIC_VECTOR'("000000"), (memory_1_mux1h_5_nl
      & memory_1_mux1h_12_nl & memory_1_mux1h_13_nl), memory_1_nor_1_seb);
  memory_1_mux1h_6_nl <= MUX1HOT_s_1_7_2((z_out_12(0)), (z_out_4(0)), (z_out_23(0)),
      (z_out_25(0)), (z_out_20(1)), (z_out_21(1)), (perceptron_simple_k_7_0_sva(3)),
      STD_LOGIC_VECTOR'( memory_1_or_2_cse & and_316_cse & memory_1_or_5_cse & and_318_cse
      & memory_1_or_6_cse_1 & and_317_cse & (fsm_output(87))));
  memory_1_and_5_nl <= memory_1_mux1h_6_nl AND memory_1_nor_1_seb;
  memory_1_mux1h_7_nl <= MUX1HOT_s_1_8_2((CR1_simple_j_2_4_0_sva(2)), (CR1_simple_j_4_0_sva(2)),
      (FOR_A_1_oelse_acc_1_ncse_sva_2(1)), (z_out_8(0)), (z_out_4(0)), (z_out_20(0)),
      (z_out_21(0)), (perceptron_simple_k_7_0_sva(2)), STD_LOGIC_VECTOR'( (fsm_output(10))
      & (fsm_output(15)) & and_316_cse & memory_1_or_5_cse & and_318_cse & memory_1_or_6_cse_1
      & and_317_cse & (fsm_output(87))));
  memory_1_and_6_nl <= memory_1_mux1h_7_nl AND memory_1_nor_1_seb;
  memory_1_mux1h_8_nl <= MUX1HOT_s_1_9_2((CR1_simple_j_2_4_0_sva(1)), (CR1_simple_j_4_0_sva(1)),
      (FOR_A_1_oelse_acc_1_ncse_sva_2(0)), (CR2_simple_j_2_3_0_sva(1)), (CR2_simple_j_3_0_sva(1)),
      (FOR_A_3_oelse_acc_1_ncse_sva_2(0)), (z_out_27_2_0(0)), (z_out_4(0)), (perceptron_simple_k_7_0_sva(1)),
      STD_LOGIC_VECTOR'( (fsm_output(10)) & (fsm_output(15)) & and_316_cse & (fsm_output(36))
      & (fsm_output(41)) & and_318_cse & memory_1_or_6_cse_1 & and_317_cse & (fsm_output(87))));
  memory_1_and_7_nl <= memory_1_mux1h_8_nl AND memory_1_nor_1_seb;
  memory_1_mux1h_9_nl <= MUX1HOT_s_1_10_2((CR1_simple_j_2_4_0_sva(0)), (CR1_simple_j_4_0_sva(0)),
      (MP1_simple_a_1_0_sva(0)), (CR2_simple_j_2_3_0_sva(0)), (CR2_simple_j_3_0_sva(0)),
      (MP2_simple_a_1_0_sva(0)), (CR3_simple_j_2_2_0_sva(0)), (CR3_simple_j_2_0_sva(0)),
      (MP3_simple_a_1_0_sva(0)), (perceptron_simple_k_7_0_sva(0)), STD_LOGIC_VECTOR'(
      (fsm_output(10)) & (fsm_output(15)) & and_316_cse & (fsm_output(36)) & (fsm_output(41))
      & and_318_cse & (fsm_output(62)) & (fsm_output(67)) & and_317_cse & (fsm_output(87))));
  memory_1_and_8_nl <= memory_1_mux1h_9_nl AND memory_1_nor_1_seb;
  memory_1_rsci_radr_d <= memory_1_and_1_nl & memory_1_and_4_nl & memory_1_and_5_nl
      & memory_1_and_6_nl & memory_1_and_7_nl & memory_1_and_8_nl;
  reshape_simple_add_N_or_cse <= (fsm_output(11)) OR (fsm_output(16));
  reshape_simple_add_N_or_11_cse <= (fsm_output(37)) OR (fsm_output(42));
  reshape_simple_add_N_or_2_cse <= (fsm_output(63)) OR (fsm_output(68));
  reshape_simple_add_N_mux1h_nl <= MUX1HOT_s_1_5_2((reshape_simple_add_N_10_0_lpi_4(10)),
      (INIT_I_asn_CR1_simple_add_AF_10_INIT_I_acc_sdt(4)), (reg_FOR_I_asn_CR1_simple_add_AF_10_FOR_I_acc_psp_cse(4)),
      (z_out_7(3)), (reg_FOR_I_2_acc_11_psp_cse(3)), STD_LOGIC_VECTOR'( or_220_ssc
      & (fsm_output(3)) & reshape_simple_add_N_or_cse & (fsm_output(29)) & reshape_simple_add_N_or_11_cse));
  reshape_simple_add_N_and_nl <= reshape_simple_add_N_mux1h_nl AND (NOT((fsm_output(55))
      OR (fsm_output(63)) OR (fsm_output(68)))) AND memory_1_or_1_seb;
  reshape_simple_add_N_mux1h_4_nl <= MUX1HOT_v_4_7_2((reshape_simple_add_N_10_0_lpi_4(9
      DOWNTO 6)), (INIT_I_asn_CR1_simple_add_AF_10_INIT_I_acc_sdt(3 DOWNTO 0)), (reg_FOR_I_asn_CR1_simple_add_AF_10_FOR_I_acc_psp_cse(3
      DOWNTO 0)), ((z_out_7(2 DOWNTO 0)) & (z_out_10(2))), ((reg_FOR_I_2_acc_11_psp_cse(2
      DOWNTO 0)) & (reg_FOR_I_2_acc_9_sdt_cse(2))), (z_out_12(4 DOWNTO 1)), (reg_FOR_I_4_acc_11_psp_cse(4
      DOWNTO 1)), STD_LOGIC_VECTOR'( or_220_ssc & (fsm_output(3)) & reshape_simple_add_N_or_cse
      & (fsm_output(29)) & reshape_simple_add_N_or_11_cse & (fsm_output(55)) & reshape_simple_add_N_or_2_cse));
  reshape_simple_add_N_or_3_nl <= (fsm_output(3)) OR (fsm_output(29));
  reshape_simple_add_N_or_15_nl <= reshape_simple_add_N_or_cse OR reshape_simple_add_N_or_11_cse;
  reshape_simple_add_N_mux1h_9_nl <= MUX1HOT_v_2_5_2((reshape_simple_add_N_10_0_lpi_4(5
      DOWNTO 4)), (z_out_10(1 DOWNTO 0)), (reg_FOR_I_2_acc_9_sdt_cse(1 DOWNTO 0)),
      STD_LOGIC_VECTOR'( (z_out_12(0)) & (INIT_I_2_acc_6_sdt_1(2))), STD_LOGIC_VECTOR'(
      (reg_FOR_I_4_acc_11_psp_cse(0)) & (reg_FOR_I_4_acc_9_sdt_cse(2))), STD_LOGIC_VECTOR'(
      or_220_ssc & reshape_simple_add_N_or_3_nl & reshape_simple_add_N_or_15_nl &
      (fsm_output(55)) & reshape_simple_add_N_or_2_cse));
  reshape_simple_add_N_and_2_nl <= MUX_v_6_2_2(STD_LOGIC_VECTOR'("000000"), (reshape_simple_add_N_mux1h_4_nl
      & reshape_simple_add_N_mux1h_9_nl), memory_1_or_1_seb);
  reshape_simple_add_N_mux1h_5_nl <= MUX1HOT_s_1_7_2((reshape_simple_add_N_10_0_lpi_4(3)),
      (z_out_12(0)), (reg_FOR_I_4_acc_11_psp_cse(0)), (z_out_23(0)), reg_FOR_I_2_acc_10_psp_cse,
      (INIT_I_2_acc_6_sdt_1(1)), (reg_FOR_I_4_acc_9_sdt_cse(1)), STD_LOGIC_VECTOR'(
      or_220_ssc & (fsm_output(3)) & reshape_simple_add_N_or_cse & (fsm_output(29))
      & reshape_simple_add_N_or_11_cse & (fsm_output(55)) & reshape_simple_add_N_or_2_cse));
  reshape_simple_add_N_and_3_nl <= reshape_simple_add_N_mux1h_5_nl AND memory_1_or_1_seb;
  reshape_simple_add_N_mux1h_6_nl <= MUX1HOT_s_1_8_2((reshape_simple_add_N_10_0_lpi_4(2)),
      (CR1_simple_j_1_4_0_sva(2)), (CR1_simple_j_2_4_0_sva(2)), (CR1_simple_j_4_0_sva(2)),
      (z_out_8(0)), reg_FOR_I_2_acc_8_sdt_cse, (INIT_I_2_acc_6_sdt_1(0)), (reg_FOR_I_4_acc_9_sdt_cse(0)),
      STD_LOGIC_VECTOR'( or_220_ssc & (fsm_output(3)) & (fsm_output(11)) & (fsm_output(16))
      & (fsm_output(29)) & reshape_simple_add_N_or_11_cse & (fsm_output(55)) & reshape_simple_add_N_or_2_cse));
  reshape_simple_add_N_and_4_nl <= reshape_simple_add_N_mux1h_6_nl AND memory_1_or_1_seb;
  reshape_simple_add_N_mux1h_7_nl <= MUX1HOT_s_1_9_2((reshape_simple_add_N_10_0_lpi_4(1)),
      (CR1_simple_j_1_4_0_sva(1)), (CR1_simple_j_2_4_0_sva(1)), (CR1_simple_j_4_0_sva(1)),
      (CR2_simple_j_1_3_0_sva(1)), (CR2_simple_j_2_3_0_sva(1)), (CR2_simple_j_3_0_sva(1)),
      (z_out_27_2_0(0)), reg_FOR_I_4_acc_8_sdt_2_0_cse, STD_LOGIC_VECTOR'( or_220_ssc
      & (fsm_output(3)) & (fsm_output(11)) & (fsm_output(16)) & (fsm_output(29))
      & (fsm_output(37)) & (fsm_output(42)) & (fsm_output(55)) & reshape_simple_add_N_or_2_cse));
  reshape_simple_add_N_mux1h_10_nl <= MUX1HOT_s_1_10_2((reshape_simple_add_N_10_0_lpi_4(0)),
      (CR1_simple_j_1_4_0_sva(0)), (CR1_simple_j_2_4_0_sva(0)), (CR1_simple_j_4_0_sva(0)),
      (CR2_simple_j_1_3_0_sva(0)), (CR2_simple_j_2_3_0_sva(0)), (CR2_simple_j_3_0_sva(0)),
      (CR3_simple_j_1_2_0_sva(0)), (CR3_simple_j_2_2_0_sva(0)), (CR3_simple_j_2_0_sva(0)),
      STD_LOGIC_VECTOR'( or_220_ssc & (fsm_output(3)) & (fsm_output(11)) & (fsm_output(16))
      & (fsm_output(29)) & (fsm_output(37)) & (fsm_output(42)) & (fsm_output(55))
      & (fsm_output(63)) & (fsm_output(68))));
  reshape_simple_add_N_and_5_nl <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), STD_LOGIC_VECTOR'(
      reshape_simple_add_N_mux1h_7_nl & reshape_simple_add_N_mux1h_10_nl), memory_1_or_1_seb);
  memory_1_rsci_wadr_d <= reshape_simple_add_N_and_nl & reshape_simple_add_N_and_2_nl
      & reshape_simple_add_N_and_3_nl & reshape_simple_add_N_and_4_nl & reshape_simple_add_N_and_5_nl;
  FOR_I_nor_3_cse <= NOT(MUX_v_14_2_2((z_out_22(14 DOWNTO 1)), STD_LOGIC_VECTOR'("11111111111111"),
      FOR_I_nor_2_cse));
  FOR_I_nor_4_cse <= NOT((z_out_22(0)) OR FOR_I_nor_2_cse);
  memory_1_or_17_cse <= (fsm_output(11)) OR (fsm_output(37)) OR (fsm_output(63));
  memory_1_or_19_cse <= (fsm_output(16)) OR (fsm_output(42)) OR (fsm_output(68));
  memory_1_memory_1_mux_nl <= MUX_s_1_2_2((z_out_22(16)), (memory_2_rsci_q_d(15)),
      fsm_output(82));
  memory_1_and_nl <= memory_1_memory_1_mux_nl AND (NOT((fsm_output(16)) OR (fsm_output(42))
      OR (fsm_output(68)))) AND memory_1_or_seb;
  FOR_I_FOR_I_nor_1_nl <= NOT(MUX_v_14_2_2(FOR_I_nor_3_cse, STD_LOGIC_VECTOR'("11111111111111"),
      FOR_I_and_4_cse));
  BIAS_I_BIAS_I_nor_nl <= NOT(FOR_I_nor_3_cse OR STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(FOR_I_and_4_cse,
      1),14)) OR STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(z_out_22(16), 1),14)));
  memory_1_mux1h_10_nl <= MUX1HOT_v_14_3_2(FOR_I_FOR_I_nor_1_nl, BIAS_I_BIAS_I_nor_nl,
      (memory_2_rsci_q_d(14 DOWNTO 1)), STD_LOGIC_VECTOR'( memory_1_or_17_cse & memory_1_or_19_cse
      & (fsm_output(82))));
  memory_1_and_9_nl <= MUX_v_14_2_2(STD_LOGIC_VECTOR'("00000000000000"), memory_1_mux1h_10_nl,
      memory_1_or_seb);
  FOR_I_FOR_I_nor_2_nl <= NOT(FOR_I_nor_4_cse OR FOR_I_and_4_cse);
  BIAS_I_BIAS_I_nor_3_nl <= NOT(FOR_I_nor_4_cse OR (z_out_22(16)));
  memory_1_mux1h_11_nl <= MUX1HOT_s_1_3_2(FOR_I_FOR_I_nor_2_nl, BIAS_I_BIAS_I_nor_3_nl,
      (memory_2_rsci_q_d(0)), STD_LOGIC_VECTOR'( memory_1_or_17_cse & memory_1_or_19_cse
      & (fsm_output(82))));
  memory_1_and_10_nl <= memory_1_mux1h_11_nl AND memory_1_or_seb;
  memory_1_rsci_d_d <= memory_1_and_nl & memory_1_and_9_nl & memory_1_and_10_nl;
  memory_1_rsci_we_d <= or_dcpl_53 OR (fsm_output(68)) OR (fsm_output(55)) OR (fsm_output(29))
      OR (fsm_output(3)) OR (fsm_output(63)) OR (fsm_output(42)) OR (fsm_output(37))
      OR (fsm_output(16)) OR (fsm_output(11)) OR (fsm_output(82));
  memory_1_rsci_re_d <= (fsm_output(62)) OR (fsm_output(36)) OR (fsm_output(10))
      OR (fsm_output(67)) OR (fsm_output(41)) OR (fsm_output(15)) OR (fsm_output(87))
      OR and_316_cse OR and_317_cse OR and_318_cse;
  FOR_B_2_if_acc_12_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(FOR_B_2_if_acc_8_sdt_1(6
      DOWNTO 3)) + UNSIGNED(CR2_simple_k_6_0_sva_5_0_1(3 DOWNTO 0)), 4));
  FOR_B_4_if_acc_16_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_SIGNED(SIGNED(FOR_B_4_if_acc_11_sdt_1(6
      DOWNTO 3)), 4), 6) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(CR3_simple_k_5_0_sva_4_0),
      5), 6), 6));
  memory_2_mux1h_1_nl <= MUX1HOT_v_8_3_2((STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(FOR_B_2_if_acc_12_nl),
      4)) & (FOR_B_2_if_acc_8_sdt_1(2 DOWNTO 0)) & (FOR_B_2_if_acc_9_psp_1(0))),
      (STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(FOR_B_4_if_acc_16_nl), 6)) & (FOR_B_4_if_acc_11_sdt_1(2
      DOWNTO 1))), (STD_LOGIC_VECTOR'( "000") & z_out_12), STD_LOGIC_VECTOR'( and_285_cse
      & and_283_cse & (fsm_output(81))));
  memory_2_not_4_nl <= NOT memory_2_rsci_radr_d_mx0c0;
  memory_2_and_3_nl <= MUX_v_8_2_2(STD_LOGIC_VECTOR'("00000000"), memory_2_mux1h_1_nl,
      memory_2_not_4_nl);
  memory_2_mux1h_4_nl <= MUX1HOT_s_1_3_2((z_out_16(0)), (FOR_B_4_if_acc_11_sdt_1(0)),
      (z_out_11(2)), STD_LOGIC_VECTOR'( and_285_cse & and_283_cse & (fsm_output(81))));
  memory_2_and_4_nl <= memory_2_mux1h_4_nl AND (NOT memory_2_rsci_radr_d_mx0c0);
  memory_2_mux1h_5_nl <= MUX1HOT_v_2_3_2((CR2_simple_j_aux_4_0_sva_1(1 DOWNTO 0)),
      STD_LOGIC_VECTOR'( (FOR_B_4_if_acc_6_sdt_1(0)) & (CR3_simple_j_aux_3_0_sva_1(0))),
      (z_out_11(1 DOWNTO 0)), STD_LOGIC_VECTOR'( and_285_cse & and_283_cse & (fsm_output(81))));
  memory_2_not_6_nl <= NOT memory_2_rsci_radr_d_mx0c0;
  memory_2_and_5_nl <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), memory_2_mux1h_5_nl,
      memory_2_not_6_nl);
  memory_2_rsci_radr_d <= memory_2_and_3_nl & memory_2_and_4_nl & memory_2_and_5_nl;
  FOR_B_1_if_acc_5_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(FOR_B_1_if_acc_3_sdt_1(6
      DOWNTO 3)) + UNSIGNED(MP1_simple_k_6_0_sva_5_0(3 DOWNTO 0)), 4));
  FOR_B_3_if_acc_5_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(z_out_10(5
      DOWNTO 3)), 3), 6) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(MP2_simple_k_5_0_sva_4_0),
      5), 6), 6));
  memory_2_mux1h_nl <= MUX1HOT_v_8_3_2((STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(FOR_B_1_if_acc_5_nl),
      4)) & (FOR_B_1_if_acc_3_sdt_1(2 DOWNTO 0)) & (z_out_23(0))), (STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(FOR_B_3_if_acc_5_nl),
      6)) & (z_out_10(2 DOWNTO 1))), (STD_LOGIC_VECTOR'( "000") & z_out_12), STD_LOGIC_VECTOR'(
      (fsm_output(24)) & (fsm_output(50)) & (fsm_output(76))));
  memory_2_not_1_nl <= NOT memory_2_rsci_wadr_d_mx0c0;
  memory_2_and_nl <= MUX_v_8_2_2(STD_LOGIC_VECTOR'("00000000"), memory_2_mux1h_nl,
      memory_2_not_1_nl);
  memory_2_mux1h_2_nl <= MUX1HOT_s_1_3_2((z_out_8(0)), (z_out_10(0)), (z_out_21(2)),
      STD_LOGIC_VECTOR'( (fsm_output(24)) & (fsm_output(50)) & (fsm_output(76))));
  memory_2_and_1_nl <= memory_2_mux1h_2_nl AND (NOT memory_2_rsci_wadr_d_mx0c0);
  memory_2_mux1h_3_nl <= MUX1HOT_v_2_3_2((MP1_simple_i_N_3_0_sva_1(1 DOWNTO 0)),
      STD_LOGIC_VECTOR'( (FOR_B_3_if_acc_sdt_1(0)) & (MP2_simple_i_N_2_0_sva_1(0))),
      (z_out_21(1 DOWNTO 0)), STD_LOGIC_VECTOR'( (fsm_output(24)) & (fsm_output(50))
      & (fsm_output(76))));
  memory_2_not_3_nl <= NOT memory_2_rsci_wadr_d_mx0c0;
  memory_2_and_2_nl <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), memory_2_mux1h_3_nl,
      memory_2_not_3_nl);
  memory_2_rsci_wadr_d <= memory_2_and_nl & memory_2_and_1_nl & memory_2_and_2_nl;
  or_198_nl <= (fsm_output(24)) OR (fsm_output(0));
  MP1_simple_bigger_mux1h_nl <= MUX1HOT_v_16_3_2(MP1_simple_bigger_lpi_6_dfm_1, MP2_simple_bigger_lpi_6_dfm_1,
      MP3_simple_bigger_lpi_6_dfm_1, STD_LOGIC_VECTOR'( or_198_nl & (fsm_output(50))
      & (fsm_output(76))));
  memory_2_nand_nl <= NOT(and_dcpl_6 AND (NOT (fsm_output(24))) AND (NOT (fsm_output(0))));
  memory_2_rsci_d_d <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"), MP1_simple_bigger_mux1h_nl,
      memory_2_nand_nl);
  memory_2_rsci_we_d <= or_dcpl_53 OR (fsm_output(76)) OR (fsm_output(50)) OR (fsm_output(24));
  memory_2_rsci_re_d <= and_283_cse OR (fsm_output(81)) OR and_285_cse;
  FOR_A_1_if_mux1h_4_cse <= MUX1HOT_v_4_5_2(MP1_simple_j_4_1_sva, MP1_simple_j_N_3_0_sva_1,
      CR2_simple_i_1_3_0_sva, CR2_simple_i_2_3_0_sva, CR2_simple_i_3_0_sva, STD_LOGIC_VECTOR'(
      (fsm_output(22)) & (fsm_output(24)) & (fsm_output(29)) & (fsm_output(36)) &
      (fsm_output(41))));
  INIT_I_or_6_cse <= (fsm_output(3)) OR (fsm_output(10)) OR (fsm_output(15));
  INIT_I_or_4_cse <= (fsm_output(74)) OR (fsm_output(76));
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_index_rsc_triosy_obj_ld_cse <= '0';
        Prob_9_15_sva_2 <= '0';
        Prob_9_0_sva_2 <= '0';
        Prob_9_14_1_sva_2 <= STD_LOGIC_VECTOR'( "00000000000000");
        Prob_8_15_sva_2 <= '0';
        Prob_8_0_sva_2 <= '0';
        Prob_8_14_1_sva_2 <= STD_LOGIC_VECTOR'( "00000000000000");
        Prob_1_15_sva_2 <= '0';
        Prob_1_0_sva_2 <= '0';
        Prob_1_14_1_sva_2 <= STD_LOGIC_VECTOR'( "00000000000000");
        Prob_7_15_sva_2 <= '0';
        Prob_7_0_sva_2 <= '0';
        Prob_7_14_1_sva_2 <= STD_LOGIC_VECTOR'( "00000000000000");
        Prob_2_15_sva_2 <= '0';
        Prob_2_0_sva_2 <= '0';
        Prob_2_14_1_sva_2 <= STD_LOGIC_VECTOR'( "00000000000000");
        Prob_6_15_sva_2 <= '0';
        Prob_6_0_sva_2 <= '0';
        Prob_6_14_1_sva_2 <= STD_LOGIC_VECTOR'( "00000000000000");
        Prob_3_15_sva_2 <= '0';
        Prob_3_0_sva_2 <= '0';
        Prob_3_14_1_sva_2 <= STD_LOGIC_VECTOR'( "00000000000000");
        Prob_5_15_sva_2 <= '0';
        Prob_5_0_sva_2 <= '0';
        Prob_5_14_1_sva_2 <= STD_LOGIC_VECTOR'( "00000000000000");
        Prob_4_15_sva_2 <= '0';
        Prob_4_0_sva_2 <= '0';
        Prob_4_14_1_sva_2 <= STD_LOGIC_VECTOR'( "00000000000000");
        CR1_simple_i_1_4_0_sva <= STD_LOGIC_VECTOR'( "00000");
        reg_INIT_I_slc_INIT_I_acc_2_cse <= '0';
        CR1_simple_i_1_4_0_sva_1 <= STD_LOGIC_VECTOR'( "00000");
        CR1_simple_b_1_0_sva <= STD_LOGIC_VECTOR'( "00");
        CR1_simple_b_1_0_sva_1 <= STD_LOGIC_VECTOR'( "00");
        FOR_B_lor_2_lpi_7_dfm_st <= '0';
        CR1_simple_aux_0_lpi_7_dfm <= '0';
        CR1_simple_aux_14_1_lpi_7_dfm <= STD_LOGIC_VECTOR'( "00000000000000");
        CR1_simple_aux_15_lpi_7_dfm <= '0';
        reg_FOR_I_asn_CR1_simple_add_AF_10_FOR_I_acc_psp_cse <= STD_LOGIC_VECTOR'(
            "00000");
        CR1_simple_i_4_0_sva <= STD_LOGIC_VECTOR'( "00000");
        BIAS_I_slc_15_1_itm <= STD_LOGIC_VECTOR'( "000000000000000");
        MP1_simple_j_N_3_0_sva <= STD_LOGIC_VECTOR'( "0000");
        MP1_simple_i_N_3_0_sva <= STD_LOGIC_VECTOR'( "0000");
        MP1_simple_a_1_0_sva <= STD_LOGIC_VECTOR'( "00");
        reg_FOR_A_1_lor_lpi_6_dfm_cse <= '0';
        CR2_simple_i_1_3_0_sva <= STD_LOGIC_VECTOR'( "0000");
        CR2_simple_i_1_3_0_sva_1 <= STD_LOGIC_VECTOR'( "0000");
        CR2_simple_b_1_0_sva <= STD_LOGIC_VECTOR'( "00");
        FOR_B_2_lor_2_lpi_7_dfm_st <= '0';
        CR2_simple_aux_0_lpi_7_dfm <= '0';
        CR2_simple_aux_14_1_lpi_7_dfm <= STD_LOGIC_VECTOR'( "00000000000000");
        CR2_simple_aux_15_lpi_7_dfm <= '0';
        reg_FOR_I_2_acc_11_psp_cse <= STD_LOGIC_VECTOR'( "0000");
        reg_FOR_I_2_acc_9_sdt_cse <= STD_LOGIC_VECTOR'( "000");
        reg_FOR_I_2_acc_10_psp_cse <= '0';
        reg_FOR_I_2_acc_8_sdt_cse <= '0';
        CR2_simple_i_3_0_sva <= STD_LOGIC_VECTOR'( "0000");
        BIAS_I_1_slc_15_1_itm <= STD_LOGIC_VECTOR'( "000000000000000");
        MP2_simple_j_N_2_0_sva <= STD_LOGIC_VECTOR'( "000");
        MP2_simple_i_N_2_0_sva <= STD_LOGIC_VECTOR'( "000");
        MP2_simple_a_1_0_sva <= STD_LOGIC_VECTOR'( "00");
        CR3_simple_i_1_2_0_sva <= STD_LOGIC_VECTOR'( "000");
        CR3_simple_i_1_2_0_sva_1 <= STD_LOGIC_VECTOR'( "000");
        CR3_simple_b_1_0_sva <= STD_LOGIC_VECTOR'( "00");
        FOR_B_4_lor_2_lpi_7_dfm_st <= '0';
        CR3_simple_aux_0_lpi_7_dfm <= '0';
        CR3_simple_aux_14_1_lpi_7_dfm <= STD_LOGIC_VECTOR'( "00000000000000");
        CR3_simple_aux_15_lpi_7_dfm <= '0';
        reg_FOR_I_4_acc_11_psp_cse <= STD_LOGIC_VECTOR'( "00000");
        reg_FOR_I_4_acc_9_sdt_cse <= STD_LOGIC_VECTOR'( "000");
        reg_FOR_I_4_acc_8_sdt_2_0_cse <= '0';
        CR3_simple_i_2_0_sva <= STD_LOGIC_VECTOR'( "000");
        BIAS_I_2_slc_15_1_itm <= STD_LOGIC_VECTOR'( "000000000000000");
        MP3_simple_j_N_1_0_sva_1_1 <= '0';
        MP3_simple_j_N_1_0_sva_0 <= '0';
        MP3_simple_i_N_1_0_sva_1_1 <= '0';
        MP3_simple_i_N_1_0_sva_0 <= '0';
        reshape_simple_k_4_0_sva <= STD_LOGIC_VECTOR'( "00000");
        Prob_0_sva_2_15 <= '0';
        Prob_0_sva_2_0 <= '0';
        Prob_0_sva_2_14_1 <= STD_LOGIC_VECTOR'( "00000000000000");
        perceptron_simple_k_7_0_sva <= STD_LOGIC_VECTOR'( "00000000");
        FOR_K_7_slc_FOR_K_7_acc_6_itm <= '0';
        FOR_K_7_mux_28_itm <= '0';
        FOR_K_7_mux_29_itm <= STD_LOGIC_VECTOR'( "00000000000000");
        FOR_K_7_mux_30_itm <= '0';
        perceptron_simple_k_7_0_sva_1 <= STD_LOGIC_VECTOR'( "00000000");
        k_sva <= STD_LOGIC_VECTOR'( "0000");
        max_sva_14_1 <= STD_LOGIC_VECTOR'( "00000000000000");
        max_sva_15 <= '0';
        max_sva_0 <= '0';
      ELSE
        reg_index_rsc_triosy_obj_ld_cse <= (NOT (z_out_7(3))) AND (fsm_output(90));
        Prob_9_15_sva_2 <= MUX_s_1_2_2(FOR_K_7_mux_1_nl, Prob_9_15_sva_2, or_tmp_125);
        Prob_9_0_sva_2 <= MUX_s_1_2_2(FOR_K_7_mux_2_nl, Prob_9_0_sva_2, or_tmp_125);
        Prob_9_14_1_sva_2 <= MUX1HOT_v_14_3_2(Prob_9_14_1_sva_1, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
            Prob_9_14_1_sva_2, STD_LOGIC_VECTOR'( Prob_Prob_nor_nl & Prob_and_19_nl
            & or_tmp_125));
        Prob_8_15_sva_2 <= MUX_s_1_2_2(FOR_K_7_mux_4_nl, Prob_8_15_sva_2, or_tmp_125);
        Prob_8_0_sva_2 <= MUX_s_1_2_2(FOR_K_7_mux_5_nl, Prob_8_0_sva_2, or_tmp_125);
        Prob_8_14_1_sva_2 <= MUX1HOT_v_14_3_2(Prob_8_14_1_sva_1, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
            Prob_8_14_1_sva_2, STD_LOGIC_VECTOR'( Prob_Prob_nor_1_nl & Prob_and_17_nl
            & or_tmp_125));
        Prob_1_15_sva_2 <= MUX_s_1_2_2(FOR_K_7_mux_7_nl, Prob_1_15_sva_2, or_tmp_125);
        Prob_1_0_sva_2 <= MUX_s_1_2_2(FOR_K_7_mux_8_nl, Prob_1_0_sva_2, or_tmp_125);
        Prob_1_14_1_sva_2 <= MUX1HOT_v_14_3_2(Prob_1_14_1_sva_1, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
            Prob_1_14_1_sva_2, STD_LOGIC_VECTOR'( Prob_Prob_nor_2_nl & Prob_and_15_nl
            & or_tmp_125));
        Prob_7_15_sva_2 <= MUX_s_1_2_2(FOR_K_7_mux_10_nl, Prob_7_15_sva_2, or_tmp_125);
        Prob_7_0_sva_2 <= MUX_s_1_2_2(FOR_K_7_mux_11_nl, Prob_7_0_sva_2, or_tmp_125);
        Prob_7_14_1_sva_2 <= MUX1HOT_v_14_3_2(Prob_7_14_1_sva_1, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
            Prob_7_14_1_sva_2, STD_LOGIC_VECTOR'( Prob_Prob_nor_3_nl & Prob_and_13_nl
            & or_tmp_125));
        Prob_2_15_sva_2 <= MUX_s_1_2_2(FOR_K_7_mux_13_nl, Prob_2_15_sva_2, or_tmp_125);
        Prob_2_0_sva_2 <= MUX_s_1_2_2(FOR_K_7_mux_14_nl, Prob_2_0_sva_2, or_tmp_125);
        Prob_2_14_1_sva_2 <= MUX1HOT_v_14_3_2(Prob_2_14_1_sva_1, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
            Prob_2_14_1_sva_2, STD_LOGIC_VECTOR'( Prob_Prob_nor_4_nl & Prob_and_11_nl
            & or_tmp_125));
        Prob_6_15_sva_2 <= MUX_s_1_2_2(FOR_K_7_mux_16_nl, Prob_6_15_sva_2, or_tmp_125);
        Prob_6_0_sva_2 <= MUX_s_1_2_2(FOR_K_7_mux_17_nl, Prob_6_0_sva_2, or_tmp_125);
        Prob_6_14_1_sva_2 <= MUX1HOT_v_14_3_2(Prob_6_14_1_sva_1, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
            Prob_6_14_1_sva_2, STD_LOGIC_VECTOR'( Prob_Prob_nor_5_nl & Prob_and_9_nl
            & or_tmp_125));
        Prob_3_15_sva_2 <= MUX_s_1_2_2(FOR_K_7_mux_19_nl, Prob_3_15_sva_2, or_tmp_125);
        Prob_3_0_sva_2 <= MUX_s_1_2_2(FOR_K_7_mux_20_nl, Prob_3_0_sva_2, or_tmp_125);
        Prob_3_14_1_sva_2 <= MUX1HOT_v_14_3_2(Prob_3_14_1_sva_1, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
            Prob_3_14_1_sva_2, STD_LOGIC_VECTOR'( Prob_Prob_nor_6_nl & Prob_and_7_nl
            & or_tmp_125));
        Prob_5_15_sva_2 <= MUX_s_1_2_2(FOR_K_7_mux_22_nl, Prob_5_15_sva_2, or_tmp_125);
        Prob_5_0_sva_2 <= MUX_s_1_2_2(FOR_K_7_mux_23_nl, Prob_5_0_sva_2, or_tmp_125);
        Prob_5_14_1_sva_2 <= MUX1HOT_v_14_3_2(Prob_5_14_1_sva_1, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
            Prob_5_14_1_sva_2, STD_LOGIC_VECTOR'( Prob_Prob_nor_7_nl & Prob_and_5_nl
            & or_tmp_125));
        Prob_4_15_sva_2 <= MUX_s_1_2_2(FOR_K_7_mux_25_nl, Prob_4_15_sva_2, or_tmp_125);
        Prob_4_0_sva_2 <= MUX_s_1_2_2(FOR_K_7_mux_26_nl, Prob_4_0_sva_2, or_tmp_125);
        Prob_4_14_1_sva_2 <= MUX1HOT_v_14_3_2(Prob_4_14_1_sva_1, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
            Prob_4_14_1_sva_2, STD_LOGIC_VECTOR'( Prob_Prob_nor_8_nl & Prob_and_3_nl
            & or_tmp_125));
        CR1_simple_i_1_4_0_sva <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), CR1_simple_i_1_4_0_sva_1,
            CR1_simple_i_nor_nl);
        reg_INIT_I_slc_INIT_I_acc_2_cse <= z_out(2);
        CR1_simple_i_1_4_0_sva_1 <= z_out_9;
        CR1_simple_b_1_0_sva <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), CR1_simple_b_1_0_sva_1,
            (fsm_output(8)));
        CR1_simple_b_1_0_sva_1 <= z_out_2(1 DOWNTO 0);
        FOR_B_lor_2_lpi_7_dfm_st <= or_125_cse;
        CR1_simple_aux_0_lpi_7_dfm <= MUX_s_1_2_2(CR1_simple_aux_0_lpi_7_mx1, CR1_simple_aux_0_lpi_7_dfm,
            and_4_cse);
        CR1_simple_aux_14_1_lpi_7_dfm <= MUX_v_14_2_2(CR1_simple_aux_14_1_lpi_7_mx1,
            CR1_simple_aux_14_1_lpi_7_dfm, and_4_cse);
        CR1_simple_aux_15_lpi_7_dfm <= MUX_s_1_2_2(CR1_simple_aux_15_lpi_7_mx1, CR1_simple_aux_15_lpi_7_dfm,
            and_4_cse);
        reg_FOR_I_asn_CR1_simple_add_AF_10_FOR_I_acc_psp_cse <= z_out_19;
        CR1_simple_i_4_0_sva <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), CR1_simple_i_4_0_sva_1,
            (fsm_output(17)));
        BIAS_I_slc_15_1_itm <= B_1_rsci_q_d(15 DOWNTO 1);
        MP1_simple_j_N_3_0_sva <= MUX_v_4_2_2(MP1_simple_j_N_3_0_sva_1, STD_LOGIC_VECTOR'("1111"),
            not_408_nl);
        MP1_simple_i_N_3_0_sva <= MUX_v_4_2_2(MP1_simple_i_N_3_0_sva_1, STD_LOGIC_VECTOR'("1111"),
            MP1_simple_i_N_not_nl);
        MP1_simple_a_1_0_sva <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), CR1_simple_b_1_0_sva_1,
            MP1_simple_a_nor_nl);
        reg_FOR_A_1_lor_lpi_6_dfm_cse <= nand_cse_1;
        CR2_simple_i_1_3_0_sva <= MUX_v_4_2_2(STD_LOGIC_VECTOR'("0000"), CR2_simple_i_1_3_0_sva_1,
            (fsm_output(30)));
        CR2_simple_i_1_3_0_sva_1 <= z_out_5;
        CR2_simple_b_1_0_sva <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), CR1_simple_b_1_0_sva_1,
            (fsm_output(34)));
        FOR_B_2_lor_2_lpi_7_dfm_st <= FOR_B_2_if_FOR_B_2_if_or_cse;
        CR2_simple_aux_0_lpi_7_dfm <= MUX_s_1_2_2(CR2_simple_aux_0_lpi_7_mx1, CR2_simple_aux_0_lpi_7_dfm,
            and_10_cse);
        CR2_simple_aux_14_1_lpi_7_dfm <= MUX_v_14_2_2(CR2_simple_aux_14_1_lpi_7_mx1,
            CR2_simple_aux_14_1_lpi_7_dfm, and_10_cse);
        CR2_simple_aux_15_lpi_7_dfm <= MUX_s_1_2_2(CR2_simple_aux_15_lpi_7_mx1, CR2_simple_aux_15_lpi_7_dfm,
            and_10_cse);
        reg_FOR_I_2_acc_11_psp_cse <= z_out_7;
        reg_FOR_I_2_acc_9_sdt_cse <= z_out_10(2 DOWNTO 0);
        reg_FOR_I_2_acc_10_psp_cse <= z_out_23(0);
        reg_FOR_I_2_acc_8_sdt_cse <= z_out_8(0);
        CR2_simple_i_3_0_sva <= MUX_v_4_2_2(STD_LOGIC_VECTOR'("0000"), CR2_simple_i_3_0_sva_1,
            (fsm_output(43)));
        BIAS_I_1_slc_15_1_itm <= B_2_rsci_q_d(15 DOWNTO 1);
        MP2_simple_j_N_2_0_sva <= MUX_v_3_2_2(MP2_simple_j_N_2_0_sva_1, STD_LOGIC_VECTOR'("111"),
            not_404_nl);
        MP2_simple_i_N_2_0_sva <= MUX_v_3_2_2(MP2_simple_i_N_2_0_sva_1, STD_LOGIC_VECTOR'("111"),
            MP2_simple_i_N_not_nl);
        MP2_simple_a_1_0_sva <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), CR1_simple_b_1_0_sva_1,
            MP2_simple_a_nor_nl);
        CR3_simple_i_1_2_0_sva <= MUX_v_3_2_2(STD_LOGIC_VECTOR'("000"), CR3_simple_i_1_2_0_sva_1,
            (fsm_output(56)));
        CR3_simple_i_1_2_0_sva_1 <= z_out_6;
        CR3_simple_b_1_0_sva <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), CR1_simple_b_1_0_sva_1,
            (fsm_output(60)));
        FOR_B_4_lor_2_lpi_7_dfm_st <= FOR_B_4_if_FOR_B_4_if_or_cse;
        CR3_simple_aux_0_lpi_7_dfm <= MUX_s_1_2_2(CR3_simple_aux_0_lpi_7_mx1, CR3_simple_aux_0_lpi_7_dfm,
            and_16_cse);
        CR3_simple_aux_14_1_lpi_7_dfm <= MUX_v_14_2_2(CR3_simple_aux_14_1_lpi_7_mx1,
            CR3_simple_aux_14_1_lpi_7_dfm, and_16_cse);
        CR3_simple_aux_15_lpi_7_dfm <= MUX_s_1_2_2(CR3_simple_aux_15_lpi_7_mx1, CR3_simple_aux_15_lpi_7_dfm,
            and_16_cse);
        reg_FOR_I_4_acc_11_psp_cse <= z_out_12;
        reg_FOR_I_4_acc_9_sdt_cse <= z_out_20(2 DOWNTO 0);
        reg_FOR_I_4_acc_8_sdt_2_0_cse <= z_out_27_2_0(0);
        CR3_simple_i_2_0_sva <= MUX_v_3_2_2(STD_LOGIC_VECTOR'("000"), CR3_simple_i_2_0_sva_1,
            (fsm_output(69)));
        BIAS_I_2_slc_15_1_itm <= B_3_rsci_q_d(15 DOWNTO 1);
        MP3_simple_j_N_1_0_sva_1_1 <= NOT (fsm_output(79));
        MP3_simple_j_N_1_0_sva_0 <= (MP3_simple_j_N_1_0_sva_1(0)) OR (NOT (fsm_output(79)));
        MP3_simple_i_N_1_0_sva_1_1 <= NOT (fsm_output(78));
        MP3_simple_i_N_1_0_sva_0 <= (MP3_simple_i_N_1_0_sva_1(0)) OR (NOT (fsm_output(78)));
        reshape_simple_k_4_0_sva <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), reshape_simple_k_4_0_sva_1,
            (fsm_output(83)));
        Prob_0_sva_2_15 <= MUX_s_1_2_2(FOR_K_7_mux_28_nl, Prob_0_sva_2_15, or_tmp_376);
        Prob_0_sva_2_0 <= MUX_s_1_2_2(FOR_K_7_mux_29_nl, Prob_0_sva_2_0, or_tmp_376);
        Prob_0_sva_2_14_1 <= MUX1HOT_v_14_3_2(Prob_0_sva_1_14_1, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
            Prob_0_sva_2_14_1, STD_LOGIC_VECTOR'( Prob_Prob_nor_9_nl & Prob_and_1_nl
            & or_tmp_376));
        perceptron_simple_k_7_0_sva <= MUX_v_8_2_2(STD_LOGIC_VECTOR'("00000000"),
            perceptron_simple_k_7_0_sva_1, (fsm_output(88)));
        FOR_K_7_slc_FOR_K_7_acc_6_itm <= READSLICE_1_7(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(FOR_K_7_acc_nl),
            7)), 6);
        FOR_K_7_mux_28_itm <= MUX_s_1_10_2(Prob_0_sva_1_15, Prob_1_15_sva_1, Prob_2_15_sva_1,
            Prob_3_15_sva_1, Prob_4_15_sva_1, Prob_5_15_sva_1, Prob_6_15_sva_1, Prob_7_15_sva_1,
            Prob_8_15_sva_1, Prob_9_15_sva_1, perceptron_simple_j_3_0_sva);
        FOR_K_7_mux_29_itm <= MUX_v_14_10_2(Prob_0_sva_1_14_1, Prob_1_14_1_sva_1,
            Prob_2_14_1_sva_1, Prob_3_14_1_sva_1, Prob_4_14_1_sva_1, Prob_5_14_1_sva_1,
            Prob_6_14_1_sva_1, Prob_7_14_1_sva_1, Prob_8_14_1_sva_1, Prob_9_14_1_sva_1,
            perceptron_simple_j_3_0_sva);
        FOR_K_7_mux_30_itm <= MUX_s_1_10_2(Prob_0_sva_1_0, Prob_1_0_sva_1, Prob_2_0_sva_1,
            Prob_3_0_sva_1, Prob_4_0_sva_1, Prob_5_0_sva_1, Prob_6_0_sva_1, Prob_7_0_sva_1,
            Prob_8_0_sva_1, Prob_9_0_sva_1, perceptron_simple_j_3_0_sva);
        perceptron_simple_k_7_0_sva_1 <= perceptron_simple_k_7_0_sva_2;
        k_sva <= MUX_v_4_2_2(STD_LOGIC_VECTOR'("0000"), z_out_5, (fsm_output(90)));
        max_sva_14_1 <= MUX_v_14_2_2(Prob_0_sva_2_14_1, max_sva_14_1_mx1, fsm_output(90));
        max_sva_15 <= MUX_s_1_2_2(Prob_0_sva_2_15, for_mux_1_nl, fsm_output(90));
        max_sva_0 <= MUX_s_1_2_2(Prob_0_sva_2_0, for_mux_2_nl, fsm_output(90));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        index_rsci_idat <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (NOT((NOT (fsm_output(90))) OR (z_out_7(3)))) = '1' ) THEN
        index_rsci_idat <= max_sva_14_1_mx1(10 DOWNTO 7);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR1_simple_l_1_6_0_sva_5_0 <= STD_LOGIC_VECTOR'( "000000");
      ELSIF ( reg_CR1_simple_l_1_6_0_sva_5_CR1_simple_l_or_cse = '1' ) THEN
        CR1_simple_l_1_6_0_sva_5_0 <= MUX_v_6_2_2(STD_LOGIC_VECTOR'("000000"), (z_out_13(5
            DOWNTO 0)), CR1_simple_l_not_1_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR1_simple_j_1_4_0_sva <= STD_LOGIC_VECTOR'( "00000");
      ELSIF ( ((fsm_output(5)) OR reg_CR1_simple_l_1_6_0_sva_5_CR1_simple_l_or_cse)
          = '1' ) THEN
        CR1_simple_j_1_4_0_sva <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), z_out_9,
            CR1_simple_j_not_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR1_simple_k_1_0_sva <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( ((fsm_output(19)) OR (fsm_output(6)) OR (fsm_output(14))) = '1' ) THEN
        CR1_simple_k_1_0_sva <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), (z_out_2(1 DOWNTO
            0)), (fsm_output(14)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR1_simple_a_1_0_sva <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( (or_332_cse OR (fsm_output(9))) = '1' ) THEN
        CR1_simple_a_1_0_sva <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), (z_out_2(1 DOWNTO
            0)), (fsm_output(9)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR1_simple_l_6_0_sva_5_0_1 <= STD_LOGIC_VECTOR'( "000000");
      ELSIF ( ((fsm_output(6)) OR (fsm_output(19))) = '1' ) THEN
        CR1_simple_l_6_0_sva_5_0_1 <= MUX_v_6_2_2(STD_LOGIC_VECTOR'("000000"), (z_out_13(5
            DOWNTO 0)), (fsm_output(19)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR1_simple_aux_15_lpi_7 <= '0';
        CR1_simple_aux_14_1_lpi_7 <= STD_LOGIC_VECTOR'( "00000000000000");
        CR1_simple_aux_0_lpi_7 <= '0';
      ELSIF ( reg_CR1_simple_CR1_simple_aux_or_1_cse = '1' ) THEN
        CR1_simple_aux_15_lpi_7 <= CR1_simple_aux_mux_14_nl AND (NOT or_332_cse);
        CR1_simple_aux_14_1_lpi_7 <= MUX_v_14_2_2(STD_LOGIC_VECTOR'("00000000000000"),
            CR1_simple_aux_mux_13_nl, not_410_nl);
        CR1_simple_aux_0_lpi_7 <= CR1_simple_aux_mux_12_nl AND (NOT or_332_cse);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR1_simple_j_2_4_0_sva <= STD_LOGIC_VECTOR'( "00000");
      ELSIF ( ((fsm_output(19)) OR (fsm_output(14)) OR (fsm_output(6)) OR (fsm_output(13)))
          = '1' ) THEN
        CR1_simple_j_2_4_0_sva <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), z_out_9,
            (fsm_output(13)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR1_simple_i_2_4_0_sva <= STD_LOGIC_VECTOR'( "00000");
      ELSIF ( or_332_cse = '1' ) THEN
        CR1_simple_i_2_4_0_sva <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), CR1_simple_i_2_4_0_sva_1,
            (fsm_output(12)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        FOR_I_slc_FOR_I_acc_2_itm <= '0';
      ELSIF ( (fsm_output(10)) = '1' ) THEN
        FOR_I_slc_FOR_I_acc_2_itm <= z_out(2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR1_simple_i_2_4_0_sva_1 <= STD_LOGIC_VECTOR'( "00000");
      ELSIF ( (fsm_output(10)) = '1' ) THEN
        CR1_simple_i_2_4_0_sva_1 <= z_out_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR1_simple_j_4_0_sva <= STD_LOGIC_VECTOR'( "00000");
      ELSIF ( ((fsm_output(14)) OR (fsm_output(18))) = '1' ) THEN
        CR1_simple_j_4_0_sva <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), z_out_9,
            (fsm_output(18)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        BIAS_I_slc_BIAS_I_acc_2_itm <= '0';
      ELSIF ( (fsm_output(15)) = '1' ) THEN
        BIAS_I_slc_BIAS_I_acc_2_itm <= z_out(2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR1_simple_i_4_0_sva_1 <= STD_LOGIC_VECTOR'( "00000");
      ELSIF ( (fsm_output(15)) = '1' ) THEN
        CR1_simple_i_4_0_sva_1 <= z_out_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP1_simple_k_6_0_sva_5_0 <= STD_LOGIC_VECTOR'( "000000");
      ELSIF ( ((fsm_output(19)) OR (fsm_output(28))) = '1' ) THEN
        MP1_simple_k_6_0_sva_5_0 <= MUX_v_6_2_2(STD_LOGIC_VECTOR'("000000"), (z_out_13(5
            DOWNTO 0)), (fsm_output(28)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP1_simple_j_4_1_sva <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( ((fsm_output(28)) OR (fsm_output(19)) OR (fsm_output(27))) = '1' )
          THEN
        MP1_simple_j_4_1_sva <= MUX_v_4_2_2(STD_LOGIC_VECTOR'("0000"), z_out_5, (fsm_output(27)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP1_simple_i_4_1_sva <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( ((fsm_output(20)) OR (fsm_output(26))) = '1' ) THEN
        MP1_simple_i_4_1_sva <= MUX_v_4_2_2(STD_LOGIC_VECTOR'("0000"), z_out_5, MP1_simple_i_not_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP1_simple_j_N_3_0_sva_1 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (fsm_output(20)) = '1' ) THEN
        MP1_simple_j_N_3_0_sva_1 <= z_out_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP1_simple_b_1_0_sva <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( ((fsm_output(21)) OR (fsm_output(25))) = '1' ) THEN
        MP1_simple_b_1_0_sva <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), CR1_simple_b_1_0_sva_1,
            MP1_simple_b_not_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP1_simple_bigger_lpi_6 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( ((fsm_output(21)) OR (fsm_output(23)) OR (fsm_output(25))) = '1' )
          THEN
        MP1_simple_bigger_lpi_6 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            memory_1_mux_3_nl, MP1_simple_bigger_not_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP1_simple_i_N_3_0_sva_1 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (fsm_output(21)) = '1' ) THEN
        MP1_simple_i_N_3_0_sva_1 <= z_out_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP1_simple_bigger_lpi_6_dfm_1 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(23)) = '1' ) THEN
        MP1_simple_bigger_lpi_6_dfm_1 <= MP1_simple_bigger_lpi_6_mx1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR2_simple_l_1_5_0_sva_4_0 <= STD_LOGIC_VECTOR'( "00000");
      ELSIF ( ((fsm_output(28)) OR (fsm_output(32))) = '1' ) THEN
        CR2_simple_l_1_5_0_sva_4_0 <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), (z_out_16(4
            DOWNTO 0)), (fsm_output(32)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR2_simple_j_1_3_0_sva <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( ((fsm_output(32)) OR (fsm_output(28)) OR (fsm_output(31))) = '1' )
          THEN
        CR2_simple_j_1_3_0_sva <= MUX_v_4_2_2(STD_LOGIC_VECTOR'("0000"), z_out_5,
            (fsm_output(31)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR2_simple_k_6_0_sva_5_0_1 <= STD_LOGIC_VECTOR'( "000000");
      ELSIF ( ((fsm_output(45)) OR (fsm_output(32)) OR (fsm_output(40))) = '1' )
          THEN
        CR2_simple_k_6_0_sva_5_0_1 <= MUX_v_6_2_2(STD_LOGIC_VECTOR'("000000"), (z_out_13(5
            DOWNTO 0)), (fsm_output(40)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR2_simple_a_1_0_sva <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( (or_400_cse OR (fsm_output(35))) = '1' ) THEN
        CR2_simple_a_1_0_sva <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), (z_out_2(1 DOWNTO
            0)), (fsm_output(35)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR2_simple_l_5_0_sva_4_0_1 <= STD_LOGIC_VECTOR'( "00000");
      ELSIF ( ((fsm_output(32)) OR (fsm_output(45))) = '1' ) THEN
        CR2_simple_l_5_0_sva_4_0_1 <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), (z_out_16(4
            DOWNTO 0)), (fsm_output(45)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR2_simple_aux_15_lpi_7 <= '0';
        CR2_simple_aux_14_1_lpi_7 <= STD_LOGIC_VECTOR'( "00000000000000");
        CR2_simple_aux_0_lpi_7 <= '0';
      ELSIF ( reg_CR2_simple_CR2_simple_aux_or_1_cse = '1' ) THEN
        CR2_simple_aux_15_lpi_7 <= CR1_simple_aux_mux_11_nl AND (NOT or_400_cse);
        CR2_simple_aux_14_1_lpi_7 <= MUX_v_14_2_2(STD_LOGIC_VECTOR'("00000000000000"),
            CR1_simple_aux_mux_10_nl, not_406_nl);
        CR2_simple_aux_0_lpi_7 <= CR1_simple_aux_mux_9_nl AND (NOT or_400_cse);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR2_simple_j_2_3_0_sva <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( ((fsm_output(45)) OR (fsm_output(40)) OR (fsm_output(32)) OR (fsm_output(39)))
          = '1' ) THEN
        CR2_simple_j_2_3_0_sva <= MUX_v_4_2_2(STD_LOGIC_VECTOR'("0000"), z_out_5,
            (fsm_output(39)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR2_simple_i_2_3_0_sva <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( or_400_cse = '1' ) THEN
        CR2_simple_i_2_3_0_sva <= MUX_v_4_2_2(STD_LOGIC_VECTOR'("0000"), CR2_simple_i_2_3_0_sva_1,
            (fsm_output(38)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        FOR_I_2_slc_FOR_I_2_acc_2_itm <= '0';
      ELSIF ( (fsm_output(36)) = '1' ) THEN
        FOR_I_2_slc_FOR_I_2_acc_2_itm <= z_out(2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR2_simple_i_2_3_0_sva_1 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (fsm_output(36)) = '1' ) THEN
        CR2_simple_i_2_3_0_sva_1 <= z_out_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR2_simple_j_3_0_sva <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( ((fsm_output(40)) OR (fsm_output(44))) = '1' ) THEN
        CR2_simple_j_3_0_sva <= MUX_v_4_2_2(STD_LOGIC_VECTOR'("0000"), z_out_5, (fsm_output(44)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        BIAS_I_1_slc_BIAS_I_1_acc_2_itm <= '0';
      ELSIF ( (fsm_output(41)) = '1' ) THEN
        BIAS_I_1_slc_BIAS_I_1_acc_2_itm <= z_out(2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR2_simple_i_3_0_sva_1 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (fsm_output(41)) = '1' ) THEN
        CR2_simple_i_3_0_sva_1 <= z_out_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP2_simple_k_5_0_sva_4_0 <= STD_LOGIC_VECTOR'( "00000");
      ELSIF ( ((fsm_output(45)) OR (fsm_output(54))) = '1' ) THEN
        MP2_simple_k_5_0_sva_4_0 <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), (z_out_16(4
            DOWNTO 0)), (fsm_output(54)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP2_simple_j_3_1_sva <= STD_LOGIC_VECTOR'( "000");
      ELSIF ( ((fsm_output(54)) OR (fsm_output(45)) OR (fsm_output(53))) = '1' )
          THEN
        MP2_simple_j_3_1_sva <= MUX_v_3_2_2(STD_LOGIC_VECTOR'("000"), z_out_6, (fsm_output(53)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP2_simple_i_3_1_sva <= STD_LOGIC_VECTOR'( "000");
      ELSIF ( ((fsm_output(46)) OR (fsm_output(52))) = '1' ) THEN
        MP2_simple_i_3_1_sva <= MUX_v_3_2_2(STD_LOGIC_VECTOR'("000"), z_out_6, MP2_simple_i_not_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP2_simple_j_N_2_0_sva_1 <= STD_LOGIC_VECTOR'( "000");
      ELSIF ( (fsm_output(46)) = '1' ) THEN
        MP2_simple_j_N_2_0_sva_1 <= z_out_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP2_simple_b_1_0_sva <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( ((fsm_output(47)) OR (fsm_output(51))) = '1' ) THEN
        MP2_simple_b_1_0_sva <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), CR1_simple_b_1_0_sva_1,
            MP2_simple_b_not_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP2_simple_bigger_lpi_6 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( ((fsm_output(47)) OR (fsm_output(49)) OR (fsm_output(51))) = '1' )
          THEN
        MP2_simple_bigger_lpi_6 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            memory_1_mux_4_nl, MP2_simple_bigger_not_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP2_simple_i_N_2_0_sva_1 <= STD_LOGIC_VECTOR'( "000");
      ELSIF ( (fsm_output(47)) = '1' ) THEN
        MP2_simple_i_N_2_0_sva_1 <= z_out_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP2_simple_bigger_lpi_6_dfm_1 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(49)) = '1' ) THEN
        MP2_simple_bigger_lpi_6_dfm_1 <= MP2_simple_bigger_lpi_6_mx1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR3_simple_l_1_4_0_sva <= STD_LOGIC_VECTOR'( "00000");
      ELSIF ( ((fsm_output(54)) OR (fsm_output(58))) = '1' ) THEN
        CR3_simple_l_1_4_0_sva <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), z_out_9,
            (fsm_output(58)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR3_simple_j_1_2_0_sva <= STD_LOGIC_VECTOR'( "000");
      ELSIF ( ((fsm_output(58)) OR (fsm_output(54)) OR (fsm_output(57))) = '1' )
          THEN
        CR3_simple_j_1_2_0_sva <= MUX_v_3_2_2(STD_LOGIC_VECTOR'("000"), z_out_6,
            (fsm_output(57)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR3_simple_k_5_0_sva_4_0 <= STD_LOGIC_VECTOR'( "00000");
      ELSIF ( ((fsm_output(71)) OR (fsm_output(58)) OR (fsm_output(66))) = '1' )
          THEN
        CR3_simple_k_5_0_sva_4_0 <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), (z_out_16(4
            DOWNTO 0)), (fsm_output(66)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR3_simple_a_1_0_sva <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( (or_468_cse OR (fsm_output(61))) = '1' ) THEN
        CR3_simple_a_1_0_sva <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), (z_out_2(1 DOWNTO
            0)), (fsm_output(61)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR3_simple_l_4_0_sva <= STD_LOGIC_VECTOR'( "00000");
      ELSIF ( ((fsm_output(58)) OR (fsm_output(71))) = '1' ) THEN
        CR3_simple_l_4_0_sva <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), z_out_9,
            (fsm_output(71)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR3_simple_aux_15_lpi_7 <= '0';
        CR3_simple_aux_14_1_lpi_7 <= STD_LOGIC_VECTOR'( "00000000000000");
        CR3_simple_aux_0_lpi_7 <= '0';
      ELSIF ( reg_CR3_simple_CR3_simple_aux_or_1_cse = '1' ) THEN
        CR3_simple_aux_15_lpi_7 <= CR1_simple_aux_mux_8_nl AND (NOT or_468_cse);
        CR3_simple_aux_14_1_lpi_7 <= MUX_v_14_2_2(STD_LOGIC_VECTOR'("00000000000000"),
            CR1_simple_aux_mux_7_nl, not_402_nl);
        CR3_simple_aux_0_lpi_7 <= CR1_simple_aux_mux_6_nl AND (NOT or_468_cse);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR3_simple_j_2_2_0_sva <= STD_LOGIC_VECTOR'( "000");
      ELSIF ( ((fsm_output(71)) OR (fsm_output(66)) OR (fsm_output(58)) OR (fsm_output(65)))
          = '1' ) THEN
        CR3_simple_j_2_2_0_sva <= MUX_v_3_2_2(STD_LOGIC_VECTOR'("000"), z_out_6,
            (fsm_output(65)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR3_simple_i_2_2_0_sva <= STD_LOGIC_VECTOR'( "000");
      ELSIF ( or_468_cse = '1' ) THEN
        CR3_simple_i_2_2_0_sva <= MUX_v_3_2_2(STD_LOGIC_VECTOR'("000"), CR3_simple_i_2_2_0_sva_1,
            (fsm_output(64)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        FOR_I_4_slc_FOR_I_4_acc_2_itm <= '0';
      ELSIF ( (fsm_output(62)) = '1' ) THEN
        FOR_I_4_slc_FOR_I_4_acc_2_itm <= z_out(2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR3_simple_i_2_2_0_sva_1 <= STD_LOGIC_VECTOR'( "000");
      ELSIF ( (fsm_output(62)) = '1' ) THEN
        CR3_simple_i_2_2_0_sva_1 <= z_out_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR3_simple_j_2_0_sva <= STD_LOGIC_VECTOR'( "000");
      ELSIF ( ((fsm_output(66)) OR (fsm_output(70))) = '1' ) THEN
        CR3_simple_j_2_0_sva <= MUX_v_3_2_2(STD_LOGIC_VECTOR'("000"), z_out_6, (fsm_output(70)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        BIAS_I_2_slc_BIAS_I_2_acc_2_itm <= '0';
      ELSIF ( (fsm_output(67)) = '1' ) THEN
        BIAS_I_2_slc_BIAS_I_2_acc_2_itm <= z_out(2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        CR3_simple_i_2_0_sva_1 <= STD_LOGIC_VECTOR'( "000");
      ELSIF ( (fsm_output(67)) = '1' ) THEN
        CR3_simple_i_2_0_sva_1 <= z_out_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP3_simple_k_4_0_sva <= STD_LOGIC_VECTOR'( "00000");
      ELSIF ( ((fsm_output(71)) OR (fsm_output(80))) = '1' ) THEN
        MP3_simple_k_4_0_sva <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), z_out_9,
            (fsm_output(80)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP3_simple_j_2_1_sva <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( ((fsm_output(71)) OR (fsm_output(80)) OR (fsm_output(79))) = '1' )
          THEN
        MP3_simple_j_2_1_sva <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), (z_out_2(1 DOWNTO
            0)), (fsm_output(79)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP3_simple_i_2_1_sva <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( ((fsm_output(72)) OR (fsm_output(78))) = '1' ) THEN
        MP3_simple_i_2_1_sva <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), (z_out_2(1 DOWNTO
            0)), MP3_simple_i_not_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP3_simple_j_N_1_0_sva_1 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( (fsm_output(72)) = '1' ) THEN
        MP3_simple_j_N_1_0_sva_1 <= z_out_2(1 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP3_simple_a_1_0_sva <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( ((fsm_output(75)) OR reg_MP3_simple_b_1_MP3_simple_b_or_cse) = '1'
          ) THEN
        MP3_simple_a_1_0_sva <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), CR1_simple_b_1_0_sva_1,
            MP3_simple_a_not_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP3_simple_b_1_0_sva <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( reg_MP3_simple_b_1_MP3_simple_b_or_cse = '1' ) THEN
        MP3_simple_b_1_0_sva <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), CR1_simple_b_1_0_sva_1,
            MP3_simple_b_not_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP3_simple_bigger_lpi_6 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( ((fsm_output(73)) OR (fsm_output(75)) OR (fsm_output(77))) = '1' )
          THEN
        MP3_simple_bigger_lpi_6 <= MUX_v_16_2_2(STD_LOGIC_VECTOR'("0000000000000000"),
            memory_1_mux_5_nl, MP3_simple_bigger_not_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP3_simple_i_N_1_0_sva_1 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( (fsm_output(73)) = '1' ) THEN
        MP3_simple_i_N_1_0_sva_1 <= z_out_2(1 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MP3_simple_bigger_lpi_6_dfm_1 <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(75)) = '1' ) THEN
        MP3_simple_bigger_lpi_6_dfm_1 <= MP3_simple_bigger_lpi_6_mx1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reshape_simple_i_1_0_sva <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( ((fsm_output(80)) OR (fsm_output(85))) = '1' ) THEN
        reshape_simple_i_1_0_sva <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), (z_out_2(1
            DOWNTO 0)), (fsm_output(85)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reshape_simple_j_1_0_sva <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( ((fsm_output(85)) OR (fsm_output(80)) OR (fsm_output(84))) = '1' )
          THEN
        reshape_simple_j_1_0_sva <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), (z_out_2(1
            DOWNTO 0)), (fsm_output(84)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reshape_simple_add_N_10_0_lpi_4 <= STD_LOGIC_VECTOR'( "00000000000");
      ELSIF ( ((fsm_output(80)) OR reshape_simple_add_N_10_0_lpi_4_mx0c1) = '1' )
          THEN
        reshape_simple_add_N_10_0_lpi_4 <= MUX_v_11_2_2(STD_LOGIC_VECTOR'("00000000000"),
            reshape_simple_add_N_10_0_sva_1, reshape_simple_add_N_10_0_lpi_4_mx0c1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        FOR_K_6_slc_FOR_K_6_acc_3_itm <= '0';
      ELSIF ( (fsm_output(81)) = '1' ) THEN
        FOR_K_6_slc_FOR_K_6_acc_3_itm <= z_out_7(3);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reshape_simple_k_4_0_sva_1 <= STD_LOGIC_VECTOR'( "00000");
      ELSIF ( (fsm_output(81)) = '1' ) THEN
        reshape_simple_k_4_0_sva_1 <= z_out_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reshape_simple_add_N_10_0_sva_1 <= STD_LOGIC_VECTOR'( "00000000000");
      ELSIF ( (NOT(CONV_SL_1_1(fsm_output(84 DOWNTO 82)/=STD_LOGIC_VECTOR'("000"))))
          = '1' ) THEN
        reshape_simple_add_N_10_0_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(reshape_simple_add_N_10_0_lpi_4)
            + UNSIGNED'( "00000000001"), 11));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        perceptron_simple_j_3_0_sva <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( ((fsm_output(85)) OR (fsm_output(89))) = '1' ) THEN
        perceptron_simple_j_3_0_sva <= MUX_v_4_2_2(STD_LOGIC_VECTOR'("0000"), z_out_5,
            (fsm_output(89)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_9_15_sva_1 <= '0';
      ELSIF ( FOR_J_7_or_29_rgt = '0' ) THEN
        Prob_9_15_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d(15)), Prob_9_15_sva_2, (FOR_K_7_acc_7_psp_sva_1(16)),
            STD_LOGIC_VECTOR'( or_tmp_379 & or_tmp_380 & FOR_J_7_and_81_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        FOR_J_7_and_21_cse_sva <= '0';
      ELSIF ( or_tmp_383 = '0' ) THEN
        FOR_J_7_and_21_cse_sva <= FOR_J_7_and_stg_2_1_sva_1 AND (perceptron_simple_j_3_0_sva(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_9_0_sva_1 <= '0';
      ELSIF ( FOR_J_7_or_29_rgt = '0' ) THEN
        Prob_9_0_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d(4)), Prob_9_0_sva_2, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
            STD_LOGIC_VECTOR'( or_tmp_379 & or_tmp_380 & FOR_J_7_and_81_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_9_14_1_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000");
      ELSIF ( FOR_J_7_or_29_rgt = '0' ) THEN
        Prob_9_14_1_sva_1 <= MUX1HOT_v_14_3_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(P_B_rsci_q_d(15
            DOWNTO 5)),14)), Prob_9_14_1_sva_2, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
            STD_LOGIC_VECTOR'( or_tmp_379 & or_tmp_380 & FOR_J_7_and_81_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_0_sva_1_15 <= '0';
      ELSIF ( FOR_J_7_or_2_rgt = '0' ) THEN
        Prob_0_sva_1_15 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d(15)), Prob_0_sva_2_15, (FOR_K_7_acc_7_psp_sva_1(16)),
            STD_LOGIC_VECTOR'( or_tmp_392 & or_tmp_393 & FOR_J_7_and_27_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        FOR_J_7_and_20_cse_sva <= '0';
      ELSIF ( or_tmp_383 = '0' ) THEN
        FOR_J_7_and_20_cse_sva <= FOR_J_7_and_stg_2_0_sva_1 AND (NOT (perceptron_simple_j_3_0_sva(3)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_0_sva_1_0 <= '0';
      ELSIF ( FOR_J_7_or_2_rgt = '0' ) THEN
        Prob_0_sva_1_0 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d(4)), Prob_0_sva_2_0, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
            STD_LOGIC_VECTOR'( or_tmp_392 & or_tmp_393 & FOR_J_7_and_27_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_0_sva_1_14_1 <= STD_LOGIC_VECTOR'( "00000000000000");
      ELSIF ( FOR_J_7_or_2_rgt = '0' ) THEN
        Prob_0_sva_1_14_1 <= MUX1HOT_v_14_3_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(P_B_rsci_q_d(15
            DOWNTO 5)),14)), Prob_0_sva_2_14_1, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
            STD_LOGIC_VECTOR'( or_tmp_392 & or_tmp_393 & FOR_J_7_and_27_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_8_15_sva_1 <= '0';
      ELSIF ( FOR_J_7_or_26_rgt = '0' ) THEN
        Prob_8_15_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d(15)), Prob_8_15_sva_2, (FOR_K_7_acc_7_psp_sva_1(16)),
            STD_LOGIC_VECTOR'( or_tmp_405 & or_tmp_406 & FOR_J_7_and_75_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        FOR_J_7_and_19_cse_sva <= '0';
      ELSIF ( or_tmp_383 = '0' ) THEN
        FOR_J_7_and_19_cse_sva <= FOR_J_7_and_stg_2_0_sva_1 AND (perceptron_simple_j_3_0_sva(3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_8_0_sva_1 <= '0';
      ELSIF ( FOR_J_7_or_26_rgt = '0' ) THEN
        Prob_8_0_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d(4)), Prob_8_0_sva_2, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
            STD_LOGIC_VECTOR'( or_tmp_405 & or_tmp_406 & FOR_J_7_and_75_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_8_14_1_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000");
      ELSIF ( FOR_J_7_or_26_rgt = '0' ) THEN
        Prob_8_14_1_sva_1 <= MUX1HOT_v_14_3_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(P_B_rsci_q_d(15
            DOWNTO 5)),14)), Prob_8_14_1_sva_2, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
            STD_LOGIC_VECTOR'( or_tmp_405 & or_tmp_406 & FOR_J_7_and_75_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_1_15_sva_1 <= '0';
      ELSIF ( FOR_J_7_or_23_rgt = '0' ) THEN
        Prob_1_15_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d(15)), Prob_1_15_sva_2, (FOR_K_7_acc_7_psp_sva_1(16)),
            STD_LOGIC_VECTOR'( or_tmp_418 & or_tmp_419 & FOR_J_7_and_69_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        FOR_J_7_and_18_cse_sva <= '0';
      ELSIF ( or_tmp_383 = '0' ) THEN
        FOR_J_7_and_18_cse_sva <= FOR_J_7_and_stg_2_1_sva_1 AND (NOT (perceptron_simple_j_3_0_sva(3)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_1_0_sva_1 <= '0';
      ELSIF ( FOR_J_7_or_23_rgt = '0' ) THEN
        Prob_1_0_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d(4)), Prob_1_0_sva_2, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
            STD_LOGIC_VECTOR'( or_tmp_418 & or_tmp_419 & FOR_J_7_and_69_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_1_14_1_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000");
      ELSIF ( FOR_J_7_or_23_rgt = '0' ) THEN
        Prob_1_14_1_sva_1 <= MUX1HOT_v_14_3_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(P_B_rsci_q_d(15
            DOWNTO 5)),14)), Prob_1_14_1_sva_2, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
            STD_LOGIC_VECTOR'( or_tmp_418 & or_tmp_419 & FOR_J_7_and_69_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_7_15_sva_1 <= '0';
      ELSIF ( FOR_J_7_or_20_rgt = '0' ) THEN
        Prob_7_15_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d(15)), Prob_7_15_sva_2, (FOR_K_7_acc_7_psp_sva_1(16)),
            STD_LOGIC_VECTOR'( or_tmp_431 & or_tmp_432 & FOR_J_7_and_63_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        FOR_J_7_and_17_cse_sva <= '0';
      ELSIF ( or_tmp_383 = '0' ) THEN
        FOR_J_7_and_17_cse_sva <= FOR_J_7_and_stg_1_3_sva_1 AND CONV_SL_1_1(perceptron_simple_j_3_0_sva(3
            DOWNTO 2)=STD_LOGIC_VECTOR'("01"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_7_0_sva_1 <= '0';
      ELSIF ( FOR_J_7_or_20_rgt = '0' ) THEN
        Prob_7_0_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d(4)), Prob_7_0_sva_2, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
            STD_LOGIC_VECTOR'( or_tmp_431 & or_tmp_432 & FOR_J_7_and_63_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_7_14_1_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000");
      ELSIF ( FOR_J_7_or_20_rgt = '0' ) THEN
        Prob_7_14_1_sva_1 <= MUX1HOT_v_14_3_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(P_B_rsci_q_d(15
            DOWNTO 5)),14)), Prob_7_14_1_sva_2, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
            STD_LOGIC_VECTOR'( or_tmp_431 & or_tmp_432 & FOR_J_7_and_63_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_2_15_sva_1 <= '0';
      ELSIF ( FOR_J_7_or_17_rgt = '0' ) THEN
        Prob_2_15_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d(15)), Prob_2_15_sva_2, (FOR_K_7_acc_7_psp_sva_1(16)),
            STD_LOGIC_VECTOR'( or_tmp_444 & or_tmp_445 & FOR_J_7_and_57_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        FOR_J_7_and_16_cse_sva <= '0';
      ELSIF ( or_tmp_383 = '0' ) THEN
        FOR_J_7_and_16_cse_sva <= FOR_J_7_and_stg_1_2_sva_1 AND CONV_SL_1_1(perceptron_simple_j_3_0_sva(3
            DOWNTO 2)=STD_LOGIC_VECTOR'("00"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_2_0_sva_1 <= '0';
      ELSIF ( FOR_J_7_or_17_rgt = '0' ) THEN
        Prob_2_0_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d(4)), Prob_2_0_sva_2, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
            STD_LOGIC_VECTOR'( or_tmp_444 & or_tmp_445 & FOR_J_7_and_57_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_2_14_1_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000");
      ELSIF ( FOR_J_7_or_17_rgt = '0' ) THEN
        Prob_2_14_1_sva_1 <= MUX1HOT_v_14_3_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(P_B_rsci_q_d(15
            DOWNTO 5)),14)), Prob_2_14_1_sva_2, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
            STD_LOGIC_VECTOR'( or_tmp_444 & or_tmp_445 & FOR_J_7_and_57_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_6_15_sva_1 <= '0';
      ELSIF ( FOR_J_7_or_14_rgt = '0' ) THEN
        Prob_6_15_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d(15)), Prob_6_15_sva_2, (FOR_K_7_acc_7_psp_sva_1(16)),
            STD_LOGIC_VECTOR'( or_tmp_457 & or_tmp_458 & FOR_J_7_and_51_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        FOR_J_7_and_15_cse_sva <= '0';
      ELSIF ( or_tmp_383 = '0' ) THEN
        FOR_J_7_and_15_cse_sva <= FOR_J_7_and_stg_1_2_sva_1 AND CONV_SL_1_1(perceptron_simple_j_3_0_sva(3
            DOWNTO 2)=STD_LOGIC_VECTOR'("01"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_6_0_sva_1 <= '0';
      ELSIF ( FOR_J_7_or_14_rgt = '0' ) THEN
        Prob_6_0_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d(4)), Prob_6_0_sva_2, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
            STD_LOGIC_VECTOR'( or_tmp_457 & or_tmp_458 & FOR_J_7_and_51_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_6_14_1_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000");
      ELSIF ( FOR_J_7_or_14_rgt = '0' ) THEN
        Prob_6_14_1_sva_1 <= MUX1HOT_v_14_3_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(P_B_rsci_q_d(15
            DOWNTO 5)),14)), Prob_6_14_1_sva_2, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
            STD_LOGIC_VECTOR'( or_tmp_457 & or_tmp_458 & FOR_J_7_and_51_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_3_15_sva_1 <= '0';
      ELSIF ( FOR_J_7_or_11_rgt = '0' ) THEN
        Prob_3_15_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d(15)), Prob_3_15_sva_2, (FOR_K_7_acc_7_psp_sva_1(16)),
            STD_LOGIC_VECTOR'( or_tmp_470 & or_tmp_471 & FOR_J_7_and_45_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        FOR_J_7_and_14_cse_sva <= '0';
      ELSIF ( or_tmp_383 = '0' ) THEN
        FOR_J_7_and_14_cse_sva <= FOR_J_7_and_stg_1_3_sva_1 AND CONV_SL_1_1(perceptron_simple_j_3_0_sva(3
            DOWNTO 2)=STD_LOGIC_VECTOR'("00"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_3_0_sva_1 <= '0';
      ELSIF ( FOR_J_7_or_11_rgt = '0' ) THEN
        Prob_3_0_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d(4)), Prob_3_0_sva_2, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
            STD_LOGIC_VECTOR'( or_tmp_470 & or_tmp_471 & FOR_J_7_and_45_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_3_14_1_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000");
      ELSIF ( FOR_J_7_or_11_rgt = '0' ) THEN
        Prob_3_14_1_sva_1 <= MUX1HOT_v_14_3_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(P_B_rsci_q_d(15
            DOWNTO 5)),14)), Prob_3_14_1_sva_2, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
            STD_LOGIC_VECTOR'( or_tmp_470 & or_tmp_471 & FOR_J_7_and_45_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_5_15_sva_1 <= '0';
      ELSIF ( FOR_J_7_or_8_rgt = '0' ) THEN
        Prob_5_15_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d(15)), Prob_5_15_sva_2, (FOR_K_7_acc_7_psp_sva_1(16)),
            STD_LOGIC_VECTOR'( or_tmp_483 & or_tmp_484 & FOR_J_7_and_39_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        FOR_J_7_and_13_cse_sva <= '0';
      ELSIF ( or_tmp_383 = '0' ) THEN
        FOR_J_7_and_13_cse_sva <= FOR_J_7_and_stg_1_1_sva_1 AND CONV_SL_1_1(perceptron_simple_j_3_0_sva(3
            DOWNTO 2)=STD_LOGIC_VECTOR'("01"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_5_0_sva_1 <= '0';
      ELSIF ( FOR_J_7_or_8_rgt = '0' ) THEN
        Prob_5_0_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d(4)), Prob_5_0_sva_2, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
            STD_LOGIC_VECTOR'( or_tmp_483 & or_tmp_484 & FOR_J_7_and_39_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_5_14_1_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000");
      ELSIF ( FOR_J_7_or_8_rgt = '0' ) THEN
        Prob_5_14_1_sva_1 <= MUX1HOT_v_14_3_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(P_B_rsci_q_d(15
            DOWNTO 5)),14)), Prob_5_14_1_sva_2, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
            STD_LOGIC_VECTOR'( or_tmp_483 & or_tmp_484 & FOR_J_7_and_39_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_4_15_sva_1 <= '0';
      ELSIF ( FOR_J_7_or_5_rgt = '0' ) THEN
        Prob_4_15_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d(15)), Prob_4_15_sva_2, (FOR_K_7_acc_7_psp_sva_1(16)),
            STD_LOGIC_VECTOR'( or_tmp_496 & or_tmp_497 & FOR_J_7_and_33_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        FOR_J_7_and_12_cse_sva <= '0';
      ELSIF ( or_tmp_383 = '0' ) THEN
        FOR_J_7_and_12_cse_sva <= FOR_J_7_and_stg_1_0_sva_1 AND CONV_SL_1_1(perceptron_simple_j_3_0_sva(3
            DOWNTO 2)=STD_LOGIC_VECTOR'("01"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_4_0_sva_1 <= '0';
      ELSIF ( FOR_J_7_or_5_rgt = '0' ) THEN
        Prob_4_0_sva_1 <= MUX1HOT_s_1_3_2((P_B_rsci_q_d(4)), Prob_4_0_sva_2, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
            STD_LOGIC_VECTOR'( or_tmp_496 & or_tmp_497 & FOR_J_7_and_33_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        Prob_4_14_1_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000");
      ELSIF ( FOR_J_7_or_5_rgt = '0' ) THEN
        Prob_4_14_1_sva_1 <= MUX1HOT_v_14_3_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(P_B_rsci_q_d(15
            DOWNTO 5)),14)), Prob_4_14_1_sva_2, FOR_K_7_FOR_K_7_nor_1_psp_sva_1,
            STD_LOGIC_VECTOR'( or_tmp_496 & or_tmp_497 & FOR_J_7_and_33_rgt));
      END IF;
    END IF;
  END PROCESS;
  FOR_K_7_mux_1_nl <= MUX_s_1_2_2(Prob_9_15_sva_1, (FOR_K_7_acc_7_psp_sva_1(16)),
      FOR_J_7_and_21_cse_sva);
  FOR_K_7_mux_2_nl <= MUX_s_1_2_2(Prob_9_0_sva_1, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
      FOR_J_7_and_21_cse_sva);
  Prob_Prob_nor_nl <= NOT(FOR_J_7_and_21_cse_sva OR or_tmp_125);
  Prob_and_19_nl <= FOR_J_7_and_21_cse_sva AND (NOT or_tmp_125);
  FOR_K_7_mux_4_nl <= MUX_s_1_2_2(Prob_8_15_sva_1, (FOR_K_7_acc_7_psp_sva_1(16)),
      FOR_J_7_and_19_cse_sva);
  FOR_K_7_mux_5_nl <= MUX_s_1_2_2(Prob_8_0_sva_1, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
      FOR_J_7_and_19_cse_sva);
  Prob_Prob_nor_1_nl <= NOT(FOR_J_7_and_19_cse_sva OR or_tmp_125);
  Prob_and_17_nl <= FOR_J_7_and_19_cse_sva AND (NOT or_tmp_125);
  FOR_K_7_mux_7_nl <= MUX_s_1_2_2(Prob_1_15_sva_1, (FOR_K_7_acc_7_psp_sva_1(16)),
      FOR_J_7_and_18_cse_sva);
  FOR_K_7_mux_8_nl <= MUX_s_1_2_2(Prob_1_0_sva_1, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
      FOR_J_7_and_18_cse_sva);
  Prob_Prob_nor_2_nl <= NOT(FOR_J_7_and_18_cse_sva OR or_tmp_125);
  Prob_and_15_nl <= FOR_J_7_and_18_cse_sva AND (NOT or_tmp_125);
  FOR_K_7_mux_10_nl <= MUX_s_1_2_2(Prob_7_15_sva_1, (FOR_K_7_acc_7_psp_sva_1(16)),
      FOR_J_7_and_17_cse_sva);
  FOR_K_7_mux_11_nl <= MUX_s_1_2_2(Prob_7_0_sva_1, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
      FOR_J_7_and_17_cse_sva);
  Prob_Prob_nor_3_nl <= NOT(FOR_J_7_and_17_cse_sva OR or_tmp_125);
  Prob_and_13_nl <= FOR_J_7_and_17_cse_sva AND (NOT or_tmp_125);
  FOR_K_7_mux_13_nl <= MUX_s_1_2_2(Prob_2_15_sva_1, (FOR_K_7_acc_7_psp_sva_1(16)),
      FOR_J_7_and_16_cse_sva);
  FOR_K_7_mux_14_nl <= MUX_s_1_2_2(Prob_2_0_sva_1, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
      FOR_J_7_and_16_cse_sva);
  Prob_Prob_nor_4_nl <= NOT(FOR_J_7_and_16_cse_sva OR or_tmp_125);
  Prob_and_11_nl <= FOR_J_7_and_16_cse_sva AND (NOT or_tmp_125);
  FOR_K_7_mux_16_nl <= MUX_s_1_2_2(Prob_6_15_sva_1, (FOR_K_7_acc_7_psp_sva_1(16)),
      FOR_J_7_and_15_cse_sva);
  FOR_K_7_mux_17_nl <= MUX_s_1_2_2(Prob_6_0_sva_1, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
      FOR_J_7_and_15_cse_sva);
  Prob_Prob_nor_5_nl <= NOT(FOR_J_7_and_15_cse_sva OR or_tmp_125);
  Prob_and_9_nl <= FOR_J_7_and_15_cse_sva AND (NOT or_tmp_125);
  FOR_K_7_mux_19_nl <= MUX_s_1_2_2(Prob_3_15_sva_1, (FOR_K_7_acc_7_psp_sva_1(16)),
      FOR_J_7_and_14_cse_sva);
  FOR_K_7_mux_20_nl <= MUX_s_1_2_2(Prob_3_0_sva_1, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
      FOR_J_7_and_14_cse_sva);
  Prob_Prob_nor_6_nl <= NOT(FOR_J_7_and_14_cse_sva OR or_tmp_125);
  Prob_and_7_nl <= FOR_J_7_and_14_cse_sva AND (NOT or_tmp_125);
  FOR_K_7_mux_22_nl <= MUX_s_1_2_2(Prob_5_15_sva_1, (FOR_K_7_acc_7_psp_sva_1(16)),
      FOR_J_7_and_13_cse_sva);
  FOR_K_7_mux_23_nl <= MUX_s_1_2_2(Prob_5_0_sva_1, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
      FOR_J_7_and_13_cse_sva);
  Prob_Prob_nor_7_nl <= NOT(FOR_J_7_and_13_cse_sva OR or_tmp_125);
  Prob_and_5_nl <= FOR_J_7_and_13_cse_sva AND (NOT or_tmp_125);
  FOR_K_7_mux_25_nl <= MUX_s_1_2_2(Prob_4_15_sva_1, (FOR_K_7_acc_7_psp_sva_1(16)),
      FOR_J_7_and_12_cse_sva);
  FOR_K_7_mux_26_nl <= MUX_s_1_2_2(Prob_4_0_sva_1, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
      FOR_J_7_and_12_cse_sva);
  Prob_Prob_nor_8_nl <= NOT(FOR_J_7_and_12_cse_sva OR or_tmp_125);
  Prob_and_3_nl <= FOR_J_7_and_12_cse_sva AND (NOT or_tmp_125);
  CR1_simple_i_nor_nl <= NOT((fsm_output(2)) OR (fsm_output(5)) OR (fsm_output(6)));
  not_408_nl <= NOT (fsm_output(27));
  MP1_simple_i_N_not_nl <= NOT (fsm_output(26));
  MP1_simple_a_nor_nl <= NOT((fsm_output(25)) OR (fsm_output(21)));
  not_404_nl <= NOT (fsm_output(53));
  MP2_simple_i_N_not_nl <= NOT (fsm_output(52));
  MP2_simple_a_nor_nl <= NOT((fsm_output(51)) OR (fsm_output(47)));
  FOR_K_7_mux_28_nl <= MUX_s_1_2_2(Prob_0_sva_1_15, (FOR_K_7_acc_7_psp_sva_1(16)),
      FOR_J_7_and_20_cse_sva);
  FOR_K_7_mux_29_nl <= MUX_s_1_2_2(Prob_0_sva_1_0, FOR_K_7_FOR_K_7_nor_2_psp_sva_1,
      FOR_J_7_and_20_cse_sva);
  Prob_Prob_nor_9_nl <= NOT(FOR_J_7_and_20_cse_sva OR or_tmp_376);
  Prob_and_1_nl <= FOR_J_7_and_20_cse_sva AND (NOT or_tmp_376);
  FOR_K_7_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(perceptron_simple_k_7_0_sva_2(7
      DOWNTO 2)), 6), 7) + SIGNED'( "1010011"), 7));
  for_mux_1_nl <= MUX_s_1_2_2(max_sva_15, for_slc_Prob_16_15_0_cse_sva_15_1, z_out_22(16));
  for_mux_2_nl <= MUX_s_1_2_2(max_sva_0, for_slc_Prob_16_15_0_cse_sva_0_1, z_out_22(16));
  CR1_simple_l_not_1_nl <= NOT (fsm_output(2));
  CR1_simple_j_not_nl <= NOT reg_CR1_simple_l_1_6_0_sva_5_CR1_simple_l_or_cse;
  CR1_simple_aux_mux_14_nl <= MUX_s_1_2_2(CR1_simple_aux_15_lpi_7_mx1, CR1_simple_aux_15_lpi_7_dfm,
      fsm_output(9));
  CR1_simple_aux_mux_13_nl <= MUX_v_14_2_2(CR1_simple_aux_14_1_lpi_7_mx1, CR1_simple_aux_14_1_lpi_7_dfm,
      fsm_output(9));
  not_410_nl <= NOT or_332_cse;
  CR1_simple_aux_mux_12_nl <= MUX_s_1_2_2(CR1_simple_aux_0_lpi_7_mx1, CR1_simple_aux_0_lpi_7_dfm,
      fsm_output(9));
  MP1_simple_i_not_nl <= NOT (fsm_output(20));
  MP1_simple_b_not_nl <= NOT (fsm_output(21));
  memory_1_mux_3_nl <= MUX_v_16_2_2(MP1_simple_bigger_lpi_6_mx1, MP1_simple_bigger_lpi_6_dfm_1,
      fsm_output(25));
  MP1_simple_bigger_not_nl <= NOT (fsm_output(21));
  CR1_simple_aux_mux_11_nl <= MUX_s_1_2_2(CR2_simple_aux_15_lpi_7_mx1, CR2_simple_aux_15_lpi_7_dfm,
      fsm_output(35));
  CR1_simple_aux_mux_10_nl <= MUX_v_14_2_2(CR2_simple_aux_14_1_lpi_7_mx1, CR2_simple_aux_14_1_lpi_7_dfm,
      fsm_output(35));
  not_406_nl <= NOT or_400_cse;
  CR1_simple_aux_mux_9_nl <= MUX_s_1_2_2(CR2_simple_aux_0_lpi_7_mx1, CR2_simple_aux_0_lpi_7_dfm,
      fsm_output(35));
  MP2_simple_i_not_nl <= NOT (fsm_output(46));
  MP2_simple_b_not_nl <= NOT (fsm_output(47));
  memory_1_mux_4_nl <= MUX_v_16_2_2(MP2_simple_bigger_lpi_6_mx1, MP2_simple_bigger_lpi_6_dfm_1,
      fsm_output(51));
  MP2_simple_bigger_not_nl <= NOT (fsm_output(47));
  CR1_simple_aux_mux_8_nl <= MUX_s_1_2_2(CR3_simple_aux_15_lpi_7_mx1, CR3_simple_aux_15_lpi_7_dfm,
      fsm_output(61));
  CR1_simple_aux_mux_7_nl <= MUX_v_14_2_2(CR3_simple_aux_14_1_lpi_7_mx1, CR3_simple_aux_14_1_lpi_7_dfm,
      fsm_output(61));
  not_402_nl <= NOT or_468_cse;
  CR1_simple_aux_mux_6_nl <= MUX_s_1_2_2(CR3_simple_aux_0_lpi_7_mx1, CR3_simple_aux_0_lpi_7_dfm,
      fsm_output(61));
  MP3_simple_i_not_nl <= NOT (fsm_output(72));
  MP3_simple_a_not_nl <= NOT reg_MP3_simple_b_1_MP3_simple_b_or_cse;
  MP3_simple_b_not_nl <= NOT (fsm_output(73));
  memory_1_mux_5_nl <= MUX_v_16_2_2(MP3_simple_bigger_lpi_6_mx1, MP3_simple_bigger_lpi_6_dfm_1,
      fsm_output(77));
  MP3_simple_bigger_not_nl <= NOT (fsm_output(73));
  INIT_I_or_13_nl <= (fsm_output(3)) OR (fsm_output(10)) OR (fsm_output(15)) OR (fsm_output(5))
      OR (fsm_output(13)) OR (fsm_output(18));
  INIT_I_or_14_nl <= (fsm_output(29)) OR (fsm_output(36)) OR (fsm_output(41)) OR
      (fsm_output(39)) OR (fsm_output(26)) OR (fsm_output(27)) OR (fsm_output(31))
      OR (fsm_output(44));
  INIT_I_or_15_nl <= (fsm_output(55)) OR (fsm_output(62)) OR (fsm_output(67)) OR
      (fsm_output(65)) OR (fsm_output(52)) OR (fsm_output(53)) OR (fsm_output(57))
      OR (fsm_output(70));
  INIT_I_mux1h_7_nl <= MUX1HOT_v_2_7_2((z_out_9(4 DOWNTO 3)), (z_out_5(3 DOWNTO 2)),
      (z_out_6(2 DOWNTO 1)), (NOT CR3_simple_a_1_0_sva), (FOR_A_1_oelse_acc_1_ncse_sva_2(3
      DOWNTO 2)), MP3_simple_i_2_1_sva, (FOR_A_3_oelse_acc_1_ncse_sva_2(2 DOWNTO
      1)), STD_LOGIC_VECTOR'( INIT_I_or_13_nl & INIT_I_or_14_nl & INIT_I_or_15_nl
      & (fsm_output(59)) & (fsm_output(22)) & (fsm_output(74)) & (fsm_output(48))));
  INIT_I_nor_1_nl <= NOT((fsm_output(3)) OR (fsm_output(10)) OR (fsm_output(15))
      OR (fsm_output(29)) OR (fsm_output(36)) OR (fsm_output(41)) OR (fsm_output(55))
      OR (fsm_output(62)) OR (fsm_output(67)) OR (fsm_output(59)) OR (fsm_output(5))
      OR (fsm_output(13)) OR (fsm_output(39)) OR (fsm_output(65)) OR (fsm_output(18))
      OR (fsm_output(26)) OR (fsm_output(27)) OR (fsm_output(31)) OR (fsm_output(44))
      OR (fsm_output(52)) OR (fsm_output(53)) OR (fsm_output(57)) OR (fsm_output(70))
      OR (fsm_output(22)) OR (fsm_output(48)));
  INIT_I_or_17_nl <= (fsm_output(3)) OR (fsm_output(10)) OR (fsm_output(15)) OR (fsm_output(29))
      OR (fsm_output(36)) OR (fsm_output(41)) OR (fsm_output(55)) OR (fsm_output(62))
      OR (fsm_output(67)) OR (fsm_output(5)) OR (fsm_output(13)) OR (fsm_output(39))
      OR (fsm_output(65)) OR (fsm_output(18)) OR (fsm_output(26)) OR (fsm_output(27))
      OR (fsm_output(31)) OR (fsm_output(44)) OR (fsm_output(52)) OR (fsm_output(53))
      OR (fsm_output(57)) OR (fsm_output(70)) OR (fsm_output(22)) OR (fsm_output(48));
  INIT_I_mux1h_8_nl <= MUX1HOT_v_2_3_2(STD_LOGIC_VECTOR'( "01"), CR3_simple_b_1_0_sva,
      STD_LOGIC_VECTOR'( '0' & (MP3_simple_a_1_0_sva(1))), STD_LOGIC_VECTOR'( INIT_I_or_17_nl
      & (fsm_output(59)) & (fsm_output(74))));
  acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & INIT_I_mux1h_7_nl & INIT_I_nor_1_nl)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(INIT_I_mux1h_8_nl & '1'), 3), 4), 4));
  z_out <= READSLICE_3_4(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(acc_nl), 4)), 1);
  FOR_A_3_if_acc_16_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MP2_simple_j_3_1_sva)
      + CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(MP2_simple_b_1_0_sva(1), 1), 1),
      3), 3));
  FOR_A_1_if_mux1h_9_nl <= MUX1HOT_v_2_3_2((z_out_7(3 DOWNTO 2)), (READSLICE_2_3(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(FOR_A_3_if_acc_16_nl),
      3)), 1)), MP3_simple_j_2_1_sva, STD_LOGIC_VECTOR'( (fsm_output(22)) & (fsm_output(48))
      & (fsm_output(74))));
  FOR_A_1_if_nor_3_nl <= NOT((fsm_output(22)) OR (fsm_output(48)));
  FOR_A_1_if_FOR_A_1_if_or_1_nl <= (MP3_simple_b_1_0_sva(1)) OR (fsm_output(22))
      OR (fsm_output(48));
  acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & FOR_A_1_if_mux1h_9_nl
      & FOR_A_1_if_nor_3_nl) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'( FOR_A_1_if_FOR_A_1_if_or_1_nl
      & '1'), 2), 4), 4));
  z_out_1_2 <= READSLICE_1_4(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(acc_1_nl), 4)),
      3);
  FOR_B_or_3_nl <= (fsm_output(84)) OR (fsm_output(81));
  FOR_B_mux1h_6_nl <= MUX1HOT_v_2_19_2(CR1_simple_b_1_0_sva, MP1_simple_a_1_0_sva,
      MP1_simple_b_1_0_sva, CR2_simple_b_1_0_sva, MP2_simple_a_1_0_sva, MP2_simple_b_1_0_sva,
      CR3_simple_b_1_0_sva, STD_LOGIC_VECTOR'( MP3_simple_j_N_1_0_sva_1_1 & MP3_simple_j_N_1_0_sva_0),
      STD_LOGIC_VECTOR'( MP3_simple_i_N_1_0_sva_1_1 & MP3_simple_i_N_1_0_sva_0),
      MP3_simple_a_1_0_sva, MP3_simple_b_1_0_sva, CR1_simple_k_1_0_sva, CR1_simple_a_1_0_sva,
      CR2_simple_a_1_0_sva, CR3_simple_a_1_0_sva, MP3_simple_j_2_1_sva, MP3_simple_i_2_1_sva,
      reshape_simple_i_1_0_sva, reshape_simple_j_1_0_sva, STD_LOGIC_VECTOR'( (fsm_output(7))
      & (fsm_output(22)) & (fsm_output(24)) & (fsm_output(33)) & (fsm_output(48))
      & (fsm_output(50)) & (fsm_output(59)) & (fsm_output(72)) & (fsm_output(73))
      & (fsm_output(74)) & (fsm_output(76)) & (fsm_output(14)) & (fsm_output(9))
      & (fsm_output(35)) & (fsm_output(61)) & (fsm_output(79)) & (fsm_output(78))
      & (fsm_output(85)) & FOR_B_or_3_nl));
  FOR_B_FOR_B_mux_1_nl <= MUX_v_2_2_2(STD_LOGIC_VECTOR'( "01"), reshape_simple_i_1_0_sva,
      fsm_output(81));
  z_out_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(FOR_B_mux1h_6_nl),
      3) + CONV_UNSIGNED(UNSIGNED(FOR_B_FOR_B_mux_1_nl), 3), 3));
  FOR_B_if_or_4_nl <= (fsm_output(22)) OR (fsm_output(48)) OR (fsm_output(74)) OR
      (fsm_output(76)) OR (fsm_output(33));
  FOR_B_if_mux1h_6_nl <= MUX1HOT_v_2_3_2(CR1_simple_b_1_0_sva, (z_out_4(2 DOWNTO
      1)), (z_out_2(2 DOWNTO 1)), STD_LOGIC_VECTOR'( (fsm_output(7)) & FOR_B_if_or_4_nl
      & (fsm_output(81))));
  FOR_B_if_mux1h_7_nl <= MUX1HOT_v_2_7_2(CR1_simple_a_1_0_sva, MP1_simple_b_1_0_sva,
      MP2_simple_b_1_0_sva, MP3_simple_b_1_0_sva, MP3_simple_j_N_1_0_sva_1, reshape_simple_i_1_0_sva,
      CR2_simple_a_1_0_sva, STD_LOGIC_VECTOR'( (fsm_output(7)) & (fsm_output(22))
      & (fsm_output(48)) & (fsm_output(74)) & (fsm_output(76)) & (fsm_output(81))
      & (fsm_output(33))));
  z_out_3 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(FOR_B_if_mux1h_6_nl),
      3) + CONV_UNSIGNED(UNSIGNED(FOR_B_if_mux1h_7_nl), 3), 3));
  FOR_A_1_if_mux1h_10_nl <= MUX1HOT_v_2_5_2((FOR_A_1_oelse_acc_1_ncse_sva_2(3 DOWNTO
      2)), CR2_simple_b_1_0_sva, (FOR_A_3_oelse_acc_1_ncse_sva_2(2 DOWNTO 1)), MP3_simple_i_2_1_sva,
      MP3_simple_i_N_1_0_sva_1, STD_LOGIC_VECTOR'( (fsm_output(22)) & (fsm_output(33))
      & (fsm_output(48)) & (fsm_output(74)) & (fsm_output(76))));
  FOR_A_1_if_and_1_nl <= (MP3_simple_a_1_0_sva(1)) AND (NOT((fsm_output(22)) OR (fsm_output(33))
      OR (fsm_output(48)) OR (fsm_output(76))));
  FOR_A_1_if_mux1h_11_nl <= MUX1HOT_v_2_5_2(MP1_simple_b_1_0_sva, CR2_simple_a_1_0_sva,
      MP2_simple_b_1_0_sva, MP3_simple_b_1_0_sva, MP3_simple_j_N_1_0_sva_1, STD_LOGIC_VECTOR'(
      (fsm_output(22)) & (fsm_output(33)) & (fsm_output(48)) & (fsm_output(74)) &
      (fsm_output(76))));
  acc_4_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(FOR_A_1_if_mux1h_10_nl
      & FOR_A_1_if_and_1_nl), 3), 4) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(FOR_A_1_if_mux1h_11_nl
      & '1'), 3), 4), 4));
  z_out_4 <= READSLICE_3_4(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(acc_4_nl), 4)),
      1);
  FOR_J_1_mux1h_2_nl <= MUX1HOT_v_4_12_2(MP1_simple_j_N_3_0_sva, MP1_simple_i_N_3_0_sva,
      MP1_simple_j_4_1_sva, MP1_simple_i_4_1_sva, CR2_simple_j_1_3_0_sva, CR2_simple_i_1_3_0_sva,
      CR2_simple_j_2_3_0_sva, CR2_simple_i_2_3_0_sva, CR2_simple_j_3_0_sva, CR2_simple_i_3_0_sva,
      k_sva, perceptron_simple_j_3_0_sva, STD_LOGIC_VECTOR'( (fsm_output(20)) & (fsm_output(21))
      & (fsm_output(27)) & (fsm_output(26)) & (fsm_output(31)) & (fsm_output(29))
      & (fsm_output(39)) & (fsm_output(36)) & (fsm_output(44)) & (fsm_output(41))
      & (fsm_output(90)) & (fsm_output(89))));
  z_out_5 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(FOR_J_1_mux1h_2_nl) + UNSIGNED'(
      "0001"), 4));
  FOR_J_3_mux1h_2_nl <= MUX1HOT_v_3_10_2(MP2_simple_j_N_2_0_sva, MP2_simple_i_N_2_0_sva,
      MP2_simple_j_3_1_sva, MP2_simple_i_3_1_sva, CR3_simple_j_1_2_0_sva, CR3_simple_i_1_2_0_sva,
      CR3_simple_j_2_2_0_sva, CR3_simple_i_2_2_0_sva, CR3_simple_j_2_0_sva, CR3_simple_i_2_0_sva,
      STD_LOGIC_VECTOR'( (fsm_output(46)) & (fsm_output(47)) & (fsm_output(53)) &
      (fsm_output(52)) & (fsm_output(57)) & (fsm_output(55)) & (fsm_output(65)) &
      (fsm_output(62)) & (fsm_output(70)) & (fsm_output(67))));
  z_out_6 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(FOR_J_3_mux1h_2_nl) + UNSIGNED'(
      "001"), 3));
  FOR_K_6_or_5_nl <= (fsm_output(81)) OR (fsm_output(71)) OR (fsm_output(58)) OR
      (fsm_output(80)) OR (fsm_output(90)) OR (fsm_output(89));
  FOR_K_6_mux1h_2_nl <= MUX1HOT_v_4_6_2(STD_LOGIC_VECTOR'( "1011"), ('0' & z_out_3),
      MP1_simple_j_4_1_sva, (CR2_simple_l_5_0_sva_4_0_1(3 DOWNTO 0)), (CR2_simple_l_1_5_0_sva_4_0(3
      DOWNTO 0)), (MP2_simple_k_5_0_sva_4_0(3 DOWNTO 0)), STD_LOGIC_VECTOR'( FOR_K_6_or_5_nl
      & (fsm_output(7)) & (fsm_output(22)) & memory_1_or_5_cse & (fsm_output(29))
      & (fsm_output(48))));
  or_nl <= (fsm_output(81)) OR (fsm_output(71)) OR (fsm_output(58)) OR (fsm_output(80));
  or_663_nl <= (fsm_output(29)) OR (fsm_output(36)) OR (fsm_output(41)) OR (fsm_output(48));
  mux1h_1_nl <= MUX1HOT_v_3_5_2((z_out_9(4 DOWNTO 2)), (z_out_17 & (CR1_simple_k_1_0_sva(0))),
      (STD_LOGIC_VECTOR'( "00") & (MP1_simple_b_1_0_sva(1))), (z_out_5(3 DOWNTO 1)),
      (z_out_10(5 DOWNTO 3)), STD_LOGIC_VECTOR'( or_nl & (fsm_output(7)) & (fsm_output(22))
      & or_tmp_376 & or_663_nl));
  z_out_7 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(FOR_K_6_mux1h_2_nl) + CONV_UNSIGNED(UNSIGNED(mux1h_1_nl),
      4), 4));
  FOR_A_1_if_FOR_A_1_if_and_1_nl <= (z_out_3(2)) AND (NOT((fsm_output(24)) OR (fsm_output(29))
      OR (fsm_output(36)) OR (fsm_output(41))));
  FOR_A_1_if_mux1h_12_nl <= MUX1HOT_v_2_5_2((z_out_3(1 DOWNTO 0)), (MP1_simple_i_N_3_0_sva_1(3
      DOWNTO 2)), (CR2_simple_j_1_3_0_sva(3 DOWNTO 2)), (CR2_simple_j_2_3_0_sva(3
      DOWNTO 2)), (CR2_simple_j_3_0_sva(3 DOWNTO 2)), STD_LOGIC_VECTOR'( (fsm_output(22))
      & (fsm_output(24)) & (fsm_output(29)) & (fsm_output(36)) & (fsm_output(41))));
  z_out_8 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(FOR_A_1_if_mux1h_4_cse) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(FOR_A_1_if_FOR_A_1_if_and_1_nl
      & FOR_A_1_if_mux1h_12_nl), 3), 4), 4));
  INIT_J_mux1h_2_nl <= MUX1HOT_v_5_10_2(CR1_simple_j_1_4_0_sva, CR1_simple_i_1_4_0_sva,
      CR1_simple_j_2_4_0_sva, CR1_simple_i_2_4_0_sva, CR1_simple_j_4_0_sva, CR1_simple_i_4_0_sva,
      CR3_simple_l_1_4_0_sva, CR3_simple_l_4_0_sva, MP3_simple_k_4_0_sva, reshape_simple_k_4_0_sva,
      STD_LOGIC_VECTOR'( (fsm_output(5)) & (fsm_output(3)) & (fsm_output(13)) & (fsm_output(10))
      & (fsm_output(18)) & (fsm_output(15)) & (fsm_output(58)) & (fsm_output(71))
      & (fsm_output(80)) & (fsm_output(81))));
  z_out_9 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(INIT_J_mux1h_2_nl) + UNSIGNED'(
      "00001"), 5));
  INIT_I_or_18_nl <= (fsm_output(48)) OR (fsm_output(50));
  INIT_I_mux1h_9_nl <= MUX1HOT_v_5_7_2(CR1_simple_i_1_4_0_sva, CR1_simple_i_2_4_0_sva,
      CR1_simple_i_4_0_sva, CR2_simple_l_1_5_0_sva_4_0, CR2_simple_l_5_0_sva_4_0_1,
      MP2_simple_k_5_0_sva_4_0, CR3_simple_k_5_0_sva_4_0, STD_LOGIC_VECTOR'( (fsm_output(3))
      & (fsm_output(10)) & (fsm_output(15)) & (fsm_output(29)) & memory_1_or_5_cse
      & INIT_I_or_18_nl & (fsm_output(59))));
  FOR_A_3_if_acc_17_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(z_out_25(3
      DOWNTO 1)), 3), 4) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(MP2_simple_j_3_1_sva),
      3), 4), 4));
  INIT_I_or_19_nl <= (fsm_output(29)) OR (fsm_output(36)) OR (fsm_output(41));
  INIT_I_mux1h_10_nl <= MUX1HOT_v_4_5_2((z_out_12(4 DOWNTO 1)), (z_out_23(4 DOWNTO
      1)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(FOR_A_3_if_acc_17_nl), 4)), z_out_26,
      (z_out_11(5 DOWNTO 2)), STD_LOGIC_VECTOR'( INIT_I_or_6_cse & INIT_I_or_19_nl
      & (fsm_output(48)) & (fsm_output(50)) & (fsm_output(59))));
  z_out_10 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(INIT_I_mux1h_9_nl),
      6) + CONV_UNSIGNED(UNSIGNED(INIT_I_mux1h_10_nl), 6), 6));
  FOR_B_4_if_mux_2_nl <= MUX_v_5_2_2(CR3_simple_k_5_0_sva_4_0, reshape_simple_k_4_0_sva,
      fsm_output(81));
  FOR_B_4_if_mux_3_nl <= MUX_v_4_2_2(('0' & (CR3_simple_l_4_0_sva(4 DOWNTO 2))),
      (z_out_3 & (z_out_2(0))), fsm_output(81));
  z_out_11 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(FOR_B_4_if_mux_2_nl),
      6) + CONV_UNSIGNED(UNSIGNED(FOR_B_4_if_mux_3_nl), 6), 6));
  INIT_I_mux1h_11_nl <= MUX1HOT_v_5_7_2(CR1_simple_i_1_4_0_sva, CR1_simple_i_2_4_0_sva,
      CR1_simple_i_4_0_sva, CR3_simple_l_4_0_sva, MP3_simple_k_4_0_sva, CR3_simple_l_1_4_0_sva,
      reshape_simple_k_4_0_sva, STD_LOGIC_VECTOR'( (fsm_output(3)) & (fsm_output(10))
      & (fsm_output(15)) & memory_1_or_6_cse_1 & INIT_I_or_4_cse & (fsm_output(55))
      & (fsm_output(81))));
  INIT_I_mux1h_12_nl <= MUX1HOT_v_2_7_2((CR1_simple_j_1_4_0_sva(4 DOWNTO 3)), (CR1_simple_j_2_4_0_sva(4
      DOWNTO 3)), (CR1_simple_j_4_0_sva(4 DOWNTO 3)), (z_out_20(4 DOWNTO 3)), (z_out_21(4
      DOWNTO 3)), (INIT_I_2_acc_6_sdt_1(4 DOWNTO 3)), (z_out_11(4 DOWNTO 3)), STD_LOGIC_VECTOR'(
      (fsm_output(3)) & (fsm_output(10)) & (fsm_output(15)) & memory_1_or_6_cse_1
      & INIT_I_or_4_cse & (fsm_output(55)) & (fsm_output(81))));
  z_out_12 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(INIT_I_mux1h_11_nl) + CONV_UNSIGNED(UNSIGNED(INIT_I_mux1h_12_nl),
      5), 5));
  INIT_L_mux1h_2_nl <= MUX1HOT_v_6_4_2(CR1_simple_l_1_6_0_sva_5_0, CR1_simple_l_6_0_sva_5_0_1,
      MP1_simple_k_6_0_sva_5_0, CR2_simple_k_6_0_sva_5_0_1, STD_LOGIC_VECTOR'( (fsm_output(6))
      & (fsm_output(19)) & (fsm_output(28)) & (fsm_output(40))));
  z_out_13 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(INIT_L_mux1h_2_nl),
      7) + UNSIGNED'( "0000001"), 7));
  FOR_B_mux1h_7_nl <= MUX1HOT_v_2_3_2(CR1_simple_b_1_0_sva, CR2_simple_b_1_0_sva,
      CR3_simple_a_1_0_sva, STD_LOGIC_VECTOR'( (fsm_output(7)) & (fsm_output(33))
      & (fsm_output(59))));
  z_out_14_1_0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(FOR_B_mux1h_7_nl) + UNSIGNED'(
      "11"), 2));
  FOR_B_mux1h_8_nl <= MUX1HOT_v_2_3_2(CR1_simple_a_1_0_sva, CR2_simple_a_1_0_sva,
      CR3_simple_b_1_0_sva, STD_LOGIC_VECTOR'( (fsm_output(7)) & (fsm_output(33))
      & (fsm_output(59))));
  z_out_15_1_0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(FOR_B_mux1h_8_nl) + UNSIGNED'(
      "11"), 2));
  FOR_B_mux1h_9_nl <= MUX1HOT_v_5_6_2(CR1_simple_j_2_4_0_sva, CR2_simple_l_1_5_0_sva_4_0,
      FOR_B_2_acc_1_psp_sva_1, CR2_simple_l_5_0_sva_4_0_1, MP2_simple_k_5_0_sva_4_0,
      CR3_simple_k_5_0_sva_4_0, STD_LOGIC_VECTOR'( (fsm_output(7)) & (fsm_output(32))
      & (fsm_output(33)) & (fsm_output(45)) & (fsm_output(54)) & (fsm_output(66))));
  FOR_B_or_4_nl <= (fsm_output(32)) OR (fsm_output(45)) OR (fsm_output(54)) OR (fsm_output(66));
  FOR_B_mux1h_10_nl <= MUX1HOT_v_3_3_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(z_out_14_1_0),3)),
      STD_LOGIC_VECTOR'( "001"), (CR2_simple_j_aux_4_0_sva_1(4 DOWNTO 2)), STD_LOGIC_VECTOR'(
      (fsm_output(7)) & FOR_B_or_4_nl & (fsm_output(33))));
  z_out_16 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(FOR_B_mux1h_9_nl),
      6) + CONV_UNSIGNED(SIGNED(FOR_B_mux1h_10_nl), 6), 6));
  FOR_B_if_mux1h_8_nl <= MUX1HOT_v_2_4_2(CR1_simple_b_1_0_sva, (CR1_simple_l_6_0_sva_5_0_1(1
      DOWNTO 0)), (CR1_simple_l_1_6_0_sva_5_0(1 DOWNTO 0)), (MP1_simple_k_6_0_sva_5_0(1
      DOWNTO 0)), STD_LOGIC_VECTOR'( (fsm_output(7)) & memory_1_or_2_cse & (fsm_output(3))
      & (fsm_output(22))));
  FOR_B_if_mux1h_9_nl <= MUX1HOT_s_1_3_2((CR1_simple_k_1_0_sva(1)), (z_out_10(5)),
      (z_out_23(4)), STD_LOGIC_VECTOR'( (fsm_output(7)) & INIT_I_or_6_cse & (fsm_output(22))));
  z_out_17 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(FOR_B_if_mux1h_8_nl) + CONV_UNSIGNED(CONV_UNSIGNED(FOR_B_if_mux1h_9_nl,
      1), 2), 2));
  FOR_B_if_mux1h_10_nl <= MUX1HOT_v_16_4_2(F_1_rsci_q_d, F_2_rsci_q_d, F_3_rsci_q_d,
      memory_1_rsci_q_d, STD_LOGIC_VECTOR'( (fsm_output(8)) & (fsm_output(34)) &
      (fsm_output(60)) & (fsm_output(88))));
  FOR_B_if_or_5_nl <= (fsm_output(34)) OR (fsm_output(60));
  FOR_B_if_mux1h_11_nl <= MUX1HOT_v_16_3_2(image_rsci_q_d, memory_2_rsci_q_d, P_W_rsci_q_d,
      STD_LOGIC_VECTOR'( (fsm_output(8)) & FOR_B_if_or_5_nl & (fsm_output(88))));
  mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(FOR_B_if_mux1h_10_nl)
      * SIGNED(FOR_B_if_mux1h_11_nl)), 32));
  z_out_18_31_12 <= READSLICE_20_32(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mul_nl),
      32)), 12);
  z_out_19 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(z_out_17 & (z_out_10(4 DOWNTO
      2))) + UNSIGNED(CR1_simple_l_6_0_sva_5_0_1(4 DOWNTO 0)), 5));
  z_out_20 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(CR3_simple_l_4_0_sva) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(z_out_26),
      4), 5), 5));
  FOR_A_5_if_mux_1_nl <= MUX_v_4_2_2(z_out_25, (z_out_3 & (z_out_4(0))), fsm_output(76));
  z_out_21 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MP3_simple_k_4_0_sva) + CONV_UNSIGNED(UNSIGNED(FOR_A_5_if_mux_1_nl),
      5), 5));
  FOR_I_or_3_nl <= (fsm_output(11)) OR (fsm_output(16)) OR (fsm_output(37)) OR (fsm_output(42))
      OR (fsm_output(63)) OR (fsm_output(68));
  FOR_I_mux1h_2_nl <= MUX1HOT_v_16_6_2(memory_1_rsci_q_d, MP1_simple_bigger_lpi_6,
      MP2_simple_bigger_lpi_6, ('1' & STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(NOT (CR3_simple_j_aux_3_0_sva_1(3
      DOWNTO 1))),15))), MP3_simple_bigger_lpi_6, (max_sva_15 & max_sva_14_1 & max_sva_0),
      STD_LOGIC_VECTOR'( FOR_I_or_3_nl & (fsm_output(23)) & (fsm_output(49)) & (fsm_output(59))
      & (fsm_output(75)) & (fsm_output(90))));
  FOR_I_nor_5_nl <= NOT((fsm_output(11)) OR (fsm_output(16)) OR (fsm_output(37))
      OR (fsm_output(42)) OR (fsm_output(59)) OR (fsm_output(63)) OR (fsm_output(68)));
  FOR_I_or_5_nl <= (fsm_output(23)) OR (fsm_output(49)) OR (fsm_output(75));
  FOR_I_mux1h_3_nl <= MUX1HOT_v_16_9_2((CR1_simple_aux_15_lpi_7_dfm & CR1_simple_aux_14_1_lpi_7_dfm
      & CR1_simple_aux_0_lpi_7_dfm), STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(BIAS_I_slc_15_1_itm),16)),
      (NOT memory_1_rsci_q_d), (CR2_simple_aux_15_lpi_7_dfm & CR2_simple_aux_14_1_lpi_7_dfm
      & CR2_simple_aux_0_lpi_7_dfm), STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(BIAS_I_1_slc_15_1_itm),16)),
      STD_LOGIC_VECTOR'( "0000000000000011"), (CR3_simple_aux_15_lpi_7_dfm & CR3_simple_aux_14_1_lpi_7_dfm
      & CR3_simple_aux_0_lpi_7_dfm), STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(BIAS_I_2_slc_15_1_itm),16)),
      ((NOT for_slc_Prob_16_15_0_cse_sva_15_1) & (NOT for_slc_Prob_16_15_0_cse_sva_14_1_1)
      & (NOT for_slc_Prob_16_15_0_cse_sva_0_1)), STD_LOGIC_VECTOR'( (fsm_output(11))
      & (fsm_output(16)) & FOR_I_or_5_nl & (fsm_output(37)) & (fsm_output(42)) &
      (fsm_output(59)) & (fsm_output(63)) & (fsm_output(68)) & (fsm_output(90))));
  acc_21_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_SIGNED(SIGNED(FOR_I_mux1h_2_nl
      & FOR_I_nor_5_nl), 17), 18) + CONV_UNSIGNED(CONV_SIGNED(SIGNED(FOR_I_mux1h_3_nl
      & '1'), 17), 18), 18));
  z_out_22 <= READSLICE_17_18(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(acc_21_nl),
      18)), 1);
  z_out_23 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(FOR_A_1_if_mux1h_4_cse),
      4), 5) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(z_out_8(3 DOWNTO 1)), 3), 5),
      5));
  FOR_B_2_if_mux_4_nl <= MUX_s_1_2_2(CR2_simple_aux_15_lpi_7, CR3_simple_aux_15_lpi_7,
      fsm_output(60));
  FOR_B_2_if_mux_5_nl <= MUX_v_14_2_2(CR2_simple_aux_14_1_lpi_7, CR3_simple_aux_14_1_lpi_7,
      fsm_output(60));
  FOR_B_2_if_mux_6_nl <= MUX_s_1_2_2(CR2_simple_aux_0_lpi_7, CR3_simple_aux_0_lpi_7,
      fsm_output(60));
  z_out_24 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(z_out_18_31_12) + CONV_UNSIGNED(CONV_SIGNED(SIGNED(FOR_B_2_if_mux_4_nl
      & FOR_B_2_if_mux_5_nl & FOR_B_2_if_mux_6_nl), 16), 20), 20));
  FOR_A_5_if_acc_21_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MP3_simple_j_2_1_sva)
      + CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(MP3_simple_j_2_1_sva(1), 1), 1),
      2), 2));
  FOR_A_3_if_mux_2_nl <= MUX_v_3_2_2(z_out_3, (STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(FOR_A_5_if_acc_21_nl),
      2)) & (MP3_simple_j_2_1_sva(0))), fsm_output(74));
  FOR_A_3_if_mux_3_nl <= MUX_v_3_2_2(MP2_simple_j_3_1_sva, z_out_3, fsm_output(74));
  z_out_25 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(FOR_A_3_if_mux_2_nl),
      4) + CONV_UNSIGNED(UNSIGNED(FOR_A_3_if_mux_3_nl), 4), 4));
  FOR_B_3_if_mux1h_2_nl <= MUX1HOT_v_3_4_2(MP2_simple_j_N_2_0_sva_1, CR3_simple_i_1_2_0_sva,
      CR3_simple_i_2_2_0_sva, CR3_simple_i_2_0_sva, STD_LOGIC_VECTOR'( (fsm_output(50))
      & (fsm_output(55)) & (fsm_output(62)) & (fsm_output(67))));
  FOR_B_3_if_or_1_nl <= (fsm_output(55)) OR (fsm_output(62)) OR (fsm_output(67));
  FOR_B_3_if_FOR_B_3_if_mux_1_nl <= MUX_v_2_2_2((FOR_B_3_if_acc_sdt_1(2 DOWNTO 1)),
      (z_out_27_2_0(2 DOWNTO 1)), FOR_B_3_if_or_1_nl);
  z_out_26 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(FOR_B_3_if_mux1h_2_nl),
      4) + CONV_UNSIGNED(UNSIGNED(FOR_B_3_if_FOR_B_3_if_mux_1_nl), 4), 4));
  INIT_I_2_mux1h_2_nl <= MUX1HOT_v_3_3_2(CR3_simple_i_1_2_0_sva, CR3_simple_i_2_2_0_sva,
      CR3_simple_i_2_0_sva, STD_LOGIC_VECTOR'( (fsm_output(55)) & (fsm_output(62))
      & (fsm_output(67))));
  INIT_I_2_mux1h_3_nl <= MUX1HOT_v_2_3_2((CR3_simple_j_1_2_0_sva(2 DOWNTO 1)), (CR3_simple_j_2_2_0_sva(2
      DOWNTO 1)), (CR3_simple_j_2_0_sva(2 DOWNTO 1)), STD_LOGIC_VECTOR'( (fsm_output(55))
      & (fsm_output(62)) & (fsm_output(67))));
  z_out_27_2_0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(INIT_I_2_mux1h_2_nl) +
      CONV_UNSIGNED(UNSIGNED(INIT_I_2_mux1h_3_nl), 3), 3));
END v18;

-- ------------------------------------------------------------------
--  Design Unit:    CNN_main_simple
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.BLOCK_1R1W_RBW_pkg.ALL;


ENTITY CNN_main_simple IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    image_rsc_radr : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
    image_rsc_q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    image_rsc_re : OUT STD_LOGIC;
    image_rsc_triosy_lz : OUT STD_LOGIC;
    F_1_rsc_radr : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
    F_1_rsc_q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    F_1_rsc_re : OUT STD_LOGIC;
    F_1_rsc_triosy_lz : OUT STD_LOGIC;
    B_1_rsc_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    B_1_rsc_q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    B_1_rsc_re : OUT STD_LOGIC;
    B_1_rsc_triosy_lz : OUT STD_LOGIC;
    F_2_rsc_radr : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
    F_2_rsc_q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    F_2_rsc_re : OUT STD_LOGIC;
    F_2_rsc_triosy_lz : OUT STD_LOGIC;
    B_2_rsc_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    B_2_rsc_q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    B_2_rsc_re : OUT STD_LOGIC;
    B_2_rsc_triosy_lz : OUT STD_LOGIC;
    F_3_rsc_radr : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
    F_3_rsc_q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    F_3_rsc_re : OUT STD_LOGIC;
    F_3_rsc_triosy_lz : OUT STD_LOGIC;
    B_3_rsc_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    B_3_rsc_q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    B_3_rsc_re : OUT STD_LOGIC;
    B_3_rsc_triosy_lz : OUT STD_LOGIC;
    P_W_rsc_radr : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
    P_W_rsc_q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    P_W_rsc_re : OUT STD_LOGIC;
    P_W_rsc_triosy_lz : OUT STD_LOGIC;
    P_B_rsc_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    P_B_rsc_q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    P_B_rsc_re : OUT STD_LOGIC;
    P_B_rsc_triosy_lz : OUT STD_LOGIC;
    index_rsc_dat : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    index_rsc_triosy_lz : OUT STD_LOGIC
  );
END CNN_main_simple;

ARCHITECTURE v18 OF CNN_main_simple IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL image_rsci_radr_d : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL image_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL F_1_rsci_radr_d : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL F_1_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL B_1_rsci_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL B_1_rsci_re_d : STD_LOGIC;
  SIGNAL B_1_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL F_2_rsci_radr_d : STD_LOGIC_VECTOR (14 DOWNTO 0);
  SIGNAL F_2_rsci_re_d : STD_LOGIC;
  SIGNAL F_2_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL B_2_rsci_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL B_2_rsci_re_d : STD_LOGIC;
  SIGNAL B_2_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL F_3_rsci_radr_d : STD_LOGIC_VECTOR (12 DOWNTO 0);
  SIGNAL F_3_rsci_re_d : STD_LOGIC;
  SIGNAL F_3_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL B_3_rsci_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL B_3_rsci_re_d : STD_LOGIC;
  SIGNAL B_3_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL P_W_rsci_radr_d : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL P_W_rsci_re_d : STD_LOGIC;
  SIGNAL P_W_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL P_B_rsci_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL P_B_rsci_re_d : STD_LOGIC;
  SIGNAL P_B_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL memory_1_rsci_radr_d : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL memory_1_rsci_wadr_d : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL memory_1_rsci_d_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL memory_1_rsci_we_d : STD_LOGIC;
  SIGNAL memory_1_rsci_re_d : STD_LOGIC;
  SIGNAL memory_1_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL memory_2_rsci_radr_d : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL memory_2_rsci_wadr_d : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL memory_2_rsci_d_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL memory_2_rsci_we_d : STD_LOGIC;
  SIGNAL memory_2_rsci_re_d : STD_LOGIC;
  SIGNAL memory_2_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL memory_1_rsc_we : STD_LOGIC;
  SIGNAL memory_1_rsc_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL memory_1_rsc_wadr : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL memory_1_rsc_re : STD_LOGIC;
  SIGNAL memory_1_rsc_q : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL memory_1_rsc_radr : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL memory_2_rsc_we : STD_LOGIC;
  SIGNAL memory_2_rsc_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL memory_2_rsc_wadr : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL memory_2_rsc_re : STD_LOGIC;
  SIGNAL memory_2_rsc_q : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL memory_2_rsc_radr : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL image_rsci_re_d_iff : STD_LOGIC;

  SIGNAL memory_1_rsc_comp_radr : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL memory_1_rsc_comp_wadr : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL memory_1_rsc_comp_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL memory_1_rsc_comp_q : STD_LOGIC_VECTOR (15 DOWNTO 0);

  SIGNAL memory_2_rsc_comp_radr : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL memory_2_rsc_comp_wadr : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL memory_2_rsc_comp_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL memory_2_rsc_comp_q : STD_LOGIC_VECTOR (15 DOWNTO 0);

  COMPONENT CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1728_1_gen
    PORT(
      re : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
      re_d : IN STD_LOGIC;
      q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL image_rsci_q : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL image_rsci_radr : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL image_rsci_radr_d_1 : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL image_rsci_q_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);

  COMPONENT CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1728_2_gen
    PORT(
      re : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
      re_d : IN STD_LOGIC;
      q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL F_1_rsci_q : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL F_1_rsci_radr : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL F_1_rsci_radr_d_1 : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL F_1_rsci_q_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);

  COMPONENT CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_6_64_3_gen
    PORT(
      re : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      re_d : IN STD_LOGIC;
      q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL B_1_rsci_q : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL B_1_rsci_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL B_1_rsci_radr_d_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL B_1_rsci_q_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);

  COMPONENT CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_15_18432_4_gen
    PORT(
      re : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (14 DOWNTO 0);
      re_d : IN STD_LOGIC;
      q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL F_2_rsci_q : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL F_2_rsci_radr : STD_LOGIC_VECTOR (14 DOWNTO 0);
  SIGNAL F_2_rsci_radr_d_1 : STD_LOGIC_VECTOR (14 DOWNTO 0);
  SIGNAL F_2_rsci_q_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);

  COMPONENT CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_5_32_5_gen
    PORT(
      re : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      re_d : IN STD_LOGIC;
      q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL B_2_rsci_q : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL B_2_rsci_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL B_2_rsci_radr_d_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL B_2_rsci_q_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);

  COMPONENT CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_13_5760_6_gen
    PORT(
      re : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
      re_d : IN STD_LOGIC;
      q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL F_3_rsci_q : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL F_3_rsci_radr : STD_LOGIC_VECTOR (12 DOWNTO 0);
  SIGNAL F_3_rsci_radr_d_1 : STD_LOGIC_VECTOR (12 DOWNTO 0);
  SIGNAL F_3_rsci_q_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);

  COMPONENT CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_5_20_7_gen
    PORT(
      re : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      re_d : IN STD_LOGIC;
      q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL B_3_rsci_q : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL B_3_rsci_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL B_3_rsci_radr_d_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL B_3_rsci_q_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);

  COMPONENT CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1800_8_gen
    PORT(
      re : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
      re_d : IN STD_LOGIC;
      q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL P_W_rsci_q : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL P_W_rsci_radr : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL P_W_rsci_radr_d_1 : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL P_W_rsci_q_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);

  COMPONENT CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_4_10_9_gen
    PORT(
      re : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      re_d : IN STD_LOGIC;
      q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL P_B_rsci_q : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL P_B_rsci_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL P_B_rsci_radr_d_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL P_B_rsci_q_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);

  COMPONENT CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_11_1728_11_gen
    PORT(
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
      re : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      we_d : IN STD_LOGIC;
      re_d : IN STD_LOGIC;
      q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL memory_1_rsci_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL memory_1_rsci_wadr : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL memory_1_rsci_q : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL memory_1_rsci_radr : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL memory_1_rsci_radr_d_1 : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL memory_1_rsci_wadr_d_1 : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL memory_1_rsci_d_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL memory_1_rsci_q_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);

  COMPONENT CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_11_1728_12_gen
    PORT(
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
      re : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      we_d : IN STD_LOGIC;
      re_d : IN STD_LOGIC;
      q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL memory_2_rsci_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL memory_2_rsci_wadr : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL memory_2_rsci_q : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL memory_2_rsci_radr : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL memory_2_rsci_radr_d_1 : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL memory_2_rsci_wadr_d_1 : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL memory_2_rsci_d_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL memory_2_rsci_q_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);

  COMPONENT CNN_main_simple_core
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      image_rsc_triosy_lz : OUT STD_LOGIC;
      F_1_rsc_triosy_lz : OUT STD_LOGIC;
      B_1_rsc_triosy_lz : OUT STD_LOGIC;
      F_2_rsc_triosy_lz : OUT STD_LOGIC;
      B_2_rsc_triosy_lz : OUT STD_LOGIC;
      F_3_rsc_triosy_lz : OUT STD_LOGIC;
      B_3_rsc_triosy_lz : OUT STD_LOGIC;
      P_W_rsc_triosy_lz : OUT STD_LOGIC;
      P_B_rsc_triosy_lz : OUT STD_LOGIC;
      index_rsc_dat : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      index_rsc_triosy_lz : OUT STD_LOGIC;
      image_rsci_radr_d : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
      image_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      F_1_rsci_radr_d : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
      F_1_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      B_1_rsci_radr_d : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      B_1_rsci_re_d : OUT STD_LOGIC;
      B_1_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      F_2_rsci_radr_d : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
      F_2_rsci_re_d : OUT STD_LOGIC;
      F_2_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      B_2_rsci_radr_d : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      B_2_rsci_re_d : OUT STD_LOGIC;
      B_2_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      F_3_rsci_radr_d : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
      F_3_rsci_re_d : OUT STD_LOGIC;
      F_3_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      B_3_rsci_radr_d : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      B_3_rsci_re_d : OUT STD_LOGIC;
      B_3_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      P_W_rsci_radr_d : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
      P_W_rsci_re_d : OUT STD_LOGIC;
      P_W_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      P_B_rsci_radr_d : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      P_B_rsci_re_d : OUT STD_LOGIC;
      P_B_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      memory_1_rsci_radr_d : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
      memory_1_rsci_wadr_d : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
      memory_1_rsci_d_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      memory_1_rsci_we_d : OUT STD_LOGIC;
      memory_1_rsci_re_d : OUT STD_LOGIC;
      memory_1_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      memory_2_rsci_radr_d : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
      memory_2_rsci_wadr_d : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
      memory_2_rsci_d_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      memory_2_rsci_we_d : OUT STD_LOGIC;
      memory_2_rsci_re_d : OUT STD_LOGIC;
      memory_2_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      image_rsci_re_d_pff : OUT STD_LOGIC
    );
  END COMPONENT;
  SIGNAL CNN_main_simple_core_inst_index_rsc_dat : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL CNN_main_simple_core_inst_image_rsci_radr_d : STD_LOGIC_VECTOR (10 DOWNTO
      0);
  SIGNAL CNN_main_simple_core_inst_image_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL CNN_main_simple_core_inst_F_1_rsci_radr_d : STD_LOGIC_VECTOR (10 DOWNTO
      0);
  SIGNAL CNN_main_simple_core_inst_F_1_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL CNN_main_simple_core_inst_B_1_rsci_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL CNN_main_simple_core_inst_B_1_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL CNN_main_simple_core_inst_F_2_rsci_radr_d : STD_LOGIC_VECTOR (14 DOWNTO
      0);
  SIGNAL CNN_main_simple_core_inst_F_2_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL CNN_main_simple_core_inst_B_2_rsci_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL CNN_main_simple_core_inst_B_2_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL CNN_main_simple_core_inst_F_3_rsci_radr_d : STD_LOGIC_VECTOR (12 DOWNTO
      0);
  SIGNAL CNN_main_simple_core_inst_F_3_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL CNN_main_simple_core_inst_B_3_rsci_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL CNN_main_simple_core_inst_B_3_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL CNN_main_simple_core_inst_P_W_rsci_radr_d : STD_LOGIC_VECTOR (10 DOWNTO
      0);
  SIGNAL CNN_main_simple_core_inst_P_W_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL CNN_main_simple_core_inst_P_B_rsci_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL CNN_main_simple_core_inst_P_B_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL CNN_main_simple_core_inst_memory_1_rsci_radr_d : STD_LOGIC_VECTOR (10 DOWNTO
      0);
  SIGNAL CNN_main_simple_core_inst_memory_1_rsci_wadr_d : STD_LOGIC_VECTOR (10 DOWNTO
      0);
  SIGNAL CNN_main_simple_core_inst_memory_1_rsci_d_d : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL CNN_main_simple_core_inst_memory_1_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL CNN_main_simple_core_inst_memory_2_rsci_radr_d : STD_LOGIC_VECTOR (10 DOWNTO
      0);
  SIGNAL CNN_main_simple_core_inst_memory_2_rsci_wadr_d : STD_LOGIC_VECTOR (10 DOWNTO
      0);
  SIGNAL CNN_main_simple_core_inst_memory_2_rsci_d_d : STD_LOGIC_VECTOR (15 DOWNTO
      0);
  SIGNAL CNN_main_simple_core_inst_memory_2_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO
      0);

BEGIN
  -- Default Constant Signal Assignments

  memory_1_rsc_comp : work.block_1r1w_rbw_pkg.BLOCK_1R1W_RBW
    GENERIC MAP(
      data_width => 16,
      addr_width => 11,
      depth => 1728
      )
    PORT MAP(
      radr => memory_1_rsc_comp_radr,
      wadr => memory_1_rsc_comp_wadr,
      d => memory_1_rsc_comp_d,
      we => memory_1_rsc_we,
      re => memory_1_rsc_re,
      clk => clk,
      q => memory_1_rsc_comp_q
    );
  memory_1_rsc_comp_radr <= memory_1_rsc_radr;
  memory_1_rsc_comp_wadr <= memory_1_rsc_wadr;
  memory_1_rsc_comp_d <= memory_1_rsc_d;
  memory_1_rsc_q <= memory_1_rsc_comp_q;

  memory_2_rsc_comp : work.block_1r1w_rbw_pkg.BLOCK_1R1W_RBW
    GENERIC MAP(
      data_width => 16,
      addr_width => 11,
      depth => 1728
      )
    PORT MAP(
      radr => memory_2_rsc_comp_radr,
      wadr => memory_2_rsc_comp_wadr,
      d => memory_2_rsc_comp_d,
      we => memory_2_rsc_we,
      re => memory_2_rsc_re,
      clk => clk,
      q => memory_2_rsc_comp_q
    );
  memory_2_rsc_comp_radr <= memory_2_rsc_radr;
  memory_2_rsc_comp_wadr <= memory_2_rsc_wadr;
  memory_2_rsc_comp_d <= memory_2_rsc_d;
  memory_2_rsc_q <= memory_2_rsc_comp_q;

  image_rsci : CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1728_1_gen
    PORT MAP(
      re => image_rsc_re,
      q => image_rsci_q,
      radr => image_rsci_radr,
      radr_d => image_rsci_radr_d_1,
      re_d => image_rsci_re_d_iff,
      q_d => image_rsci_q_d_1
    );
  image_rsci_q <= image_rsc_q;
  image_rsc_radr <= image_rsci_radr;
  image_rsci_radr_d_1 <= image_rsci_radr_d;
  image_rsci_q_d <= image_rsci_q_d_1;

  F_1_rsci : CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1728_2_gen
    PORT MAP(
      re => F_1_rsc_re,
      q => F_1_rsci_q,
      radr => F_1_rsci_radr,
      radr_d => F_1_rsci_radr_d_1,
      re_d => image_rsci_re_d_iff,
      q_d => F_1_rsci_q_d_1
    );
  F_1_rsci_q <= F_1_rsc_q;
  F_1_rsc_radr <= F_1_rsci_radr;
  F_1_rsci_radr_d_1 <= F_1_rsci_radr_d;
  F_1_rsci_q_d <= F_1_rsci_q_d_1;

  B_1_rsci : CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_6_64_3_gen
    PORT MAP(
      re => B_1_rsc_re,
      q => B_1_rsci_q,
      radr => B_1_rsci_radr,
      radr_d => B_1_rsci_radr_d_1,
      re_d => B_1_rsci_re_d,
      q_d => B_1_rsci_q_d_1
    );
  B_1_rsci_q <= B_1_rsc_q;
  B_1_rsc_radr <= B_1_rsci_radr;
  B_1_rsci_radr_d_1 <= B_1_rsci_radr_d;
  B_1_rsci_q_d <= B_1_rsci_q_d_1;

  F_2_rsci : CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_15_18432_4_gen
    PORT MAP(
      re => F_2_rsc_re,
      q => F_2_rsci_q,
      radr => F_2_rsci_radr,
      radr_d => F_2_rsci_radr_d_1,
      re_d => F_2_rsci_re_d,
      q_d => F_2_rsci_q_d_1
    );
  F_2_rsci_q <= F_2_rsc_q;
  F_2_rsc_radr <= F_2_rsci_radr;
  F_2_rsci_radr_d_1 <= F_2_rsci_radr_d;
  F_2_rsci_q_d <= F_2_rsci_q_d_1;

  B_2_rsci : CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_5_32_5_gen
    PORT MAP(
      re => B_2_rsc_re,
      q => B_2_rsci_q,
      radr => B_2_rsci_radr,
      radr_d => B_2_rsci_radr_d_1,
      re_d => B_2_rsci_re_d,
      q_d => B_2_rsci_q_d_1
    );
  B_2_rsci_q <= B_2_rsc_q;
  B_2_rsc_radr <= B_2_rsci_radr;
  B_2_rsci_radr_d_1 <= B_2_rsci_radr_d;
  B_2_rsci_q_d <= B_2_rsci_q_d_1;

  F_3_rsci : CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_13_5760_6_gen
    PORT MAP(
      re => F_3_rsc_re,
      q => F_3_rsci_q,
      radr => F_3_rsci_radr,
      radr_d => F_3_rsci_radr_d_1,
      re_d => F_3_rsci_re_d,
      q_d => F_3_rsci_q_d_1
    );
  F_3_rsci_q <= F_3_rsc_q;
  F_3_rsc_radr <= F_3_rsci_radr;
  F_3_rsci_radr_d_1 <= F_3_rsci_radr_d;
  F_3_rsci_q_d <= F_3_rsci_q_d_1;

  B_3_rsci : CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_5_20_7_gen
    PORT MAP(
      re => B_3_rsc_re,
      q => B_3_rsci_q,
      radr => B_3_rsci_radr,
      radr_d => B_3_rsci_radr_d_1,
      re_d => B_3_rsci_re_d,
      q_d => B_3_rsci_q_d_1
    );
  B_3_rsci_q <= B_3_rsc_q;
  B_3_rsc_radr <= B_3_rsci_radr;
  B_3_rsci_radr_d_1 <= B_3_rsci_radr_d;
  B_3_rsci_q_d <= B_3_rsci_q_d_1;

  P_W_rsci : CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_11_1800_8_gen
    PORT MAP(
      re => P_W_rsc_re,
      q => P_W_rsci_q,
      radr => P_W_rsci_radr,
      radr_d => P_W_rsci_radr_d_1,
      re_d => P_W_rsci_re_d,
      q_d => P_W_rsci_q_d_1
    );
  P_W_rsci_q <= P_W_rsc_q;
  P_W_rsc_radr <= P_W_rsci_radr;
  P_W_rsci_radr_d_1 <= P_W_rsci_radr_d;
  P_W_rsci_q_d <= P_W_rsci_q_d_1;

  P_B_rsci : CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_4_10_9_gen
    PORT MAP(
      re => P_B_rsc_re,
      q => P_B_rsci_q,
      radr => P_B_rsci_radr,
      radr_d => P_B_rsci_radr_d_1,
      re_d => P_B_rsci_re_d,
      q_d => P_B_rsci_q_d_1
    );
  P_B_rsci_q <= P_B_rsc_q;
  P_B_rsc_radr <= P_B_rsci_radr;
  P_B_rsci_radr_d_1 <= P_B_rsci_radr_d;
  P_B_rsci_q_d <= P_B_rsci_q_d_1;

  memory_1_rsci : CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_11_1728_11_gen
    PORT MAP(
      we => memory_1_rsc_we,
      d => memory_1_rsci_d,
      wadr => memory_1_rsci_wadr,
      re => memory_1_rsc_re,
      q => memory_1_rsci_q,
      radr => memory_1_rsci_radr,
      radr_d => memory_1_rsci_radr_d_1,
      wadr_d => memory_1_rsci_wadr_d_1,
      d_d => memory_1_rsci_d_d_1,
      we_d => memory_1_rsci_we_d,
      re_d => memory_1_rsci_re_d,
      q_d => memory_1_rsci_q_d_1
    );
  memory_1_rsc_d <= memory_1_rsci_d;
  memory_1_rsc_wadr <= memory_1_rsci_wadr;
  memory_1_rsci_q <= memory_1_rsc_q;
  memory_1_rsc_radr <= memory_1_rsci_radr;
  memory_1_rsci_radr_d_1 <= memory_1_rsci_radr_d;
  memory_1_rsci_wadr_d_1 <= memory_1_rsci_wadr_d;
  memory_1_rsci_d_d_1 <= memory_1_rsci_d_d;
  memory_1_rsci_q_d <= memory_1_rsci_q_d_1;

  memory_2_rsci : CNN_main_simple_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_11_1728_12_gen
    PORT MAP(
      we => memory_2_rsc_we,
      d => memory_2_rsci_d,
      wadr => memory_2_rsci_wadr,
      re => memory_2_rsc_re,
      q => memory_2_rsci_q,
      radr => memory_2_rsci_radr,
      radr_d => memory_2_rsci_radr_d_1,
      wadr_d => memory_2_rsci_wadr_d_1,
      d_d => memory_2_rsci_d_d_1,
      we_d => memory_2_rsci_we_d,
      re_d => memory_2_rsci_re_d,
      q_d => memory_2_rsci_q_d_1
    );
  memory_2_rsc_d <= memory_2_rsci_d;
  memory_2_rsc_wadr <= memory_2_rsci_wadr;
  memory_2_rsci_q <= memory_2_rsc_q;
  memory_2_rsc_radr <= memory_2_rsci_radr;
  memory_2_rsci_radr_d_1 <= memory_2_rsci_radr_d;
  memory_2_rsci_wadr_d_1 <= memory_2_rsci_wadr_d;
  memory_2_rsci_d_d_1 <= memory_2_rsci_d_d;
  memory_2_rsci_q_d <= memory_2_rsci_q_d_1;

  CNN_main_simple_core_inst : CNN_main_simple_core
    PORT MAP(
      clk => clk,
      rst => rst,
      image_rsc_triosy_lz => image_rsc_triosy_lz,
      F_1_rsc_triosy_lz => F_1_rsc_triosy_lz,
      B_1_rsc_triosy_lz => B_1_rsc_triosy_lz,
      F_2_rsc_triosy_lz => F_2_rsc_triosy_lz,
      B_2_rsc_triosy_lz => B_2_rsc_triosy_lz,
      F_3_rsc_triosy_lz => F_3_rsc_triosy_lz,
      B_3_rsc_triosy_lz => B_3_rsc_triosy_lz,
      P_W_rsc_triosy_lz => P_W_rsc_triosy_lz,
      P_B_rsc_triosy_lz => P_B_rsc_triosy_lz,
      index_rsc_dat => CNN_main_simple_core_inst_index_rsc_dat,
      index_rsc_triosy_lz => index_rsc_triosy_lz,
      image_rsci_radr_d => CNN_main_simple_core_inst_image_rsci_radr_d,
      image_rsci_q_d => CNN_main_simple_core_inst_image_rsci_q_d,
      F_1_rsci_radr_d => CNN_main_simple_core_inst_F_1_rsci_radr_d,
      F_1_rsci_q_d => CNN_main_simple_core_inst_F_1_rsci_q_d,
      B_1_rsci_radr_d => CNN_main_simple_core_inst_B_1_rsci_radr_d,
      B_1_rsci_re_d => B_1_rsci_re_d,
      B_1_rsci_q_d => CNN_main_simple_core_inst_B_1_rsci_q_d,
      F_2_rsci_radr_d => CNN_main_simple_core_inst_F_2_rsci_radr_d,
      F_2_rsci_re_d => F_2_rsci_re_d,
      F_2_rsci_q_d => CNN_main_simple_core_inst_F_2_rsci_q_d,
      B_2_rsci_radr_d => CNN_main_simple_core_inst_B_2_rsci_radr_d,
      B_2_rsci_re_d => B_2_rsci_re_d,
      B_2_rsci_q_d => CNN_main_simple_core_inst_B_2_rsci_q_d,
      F_3_rsci_radr_d => CNN_main_simple_core_inst_F_3_rsci_radr_d,
      F_3_rsci_re_d => F_3_rsci_re_d,
      F_3_rsci_q_d => CNN_main_simple_core_inst_F_3_rsci_q_d,
      B_3_rsci_radr_d => CNN_main_simple_core_inst_B_3_rsci_radr_d,
      B_3_rsci_re_d => B_3_rsci_re_d,
      B_3_rsci_q_d => CNN_main_simple_core_inst_B_3_rsci_q_d,
      P_W_rsci_radr_d => CNN_main_simple_core_inst_P_W_rsci_radr_d,
      P_W_rsci_re_d => P_W_rsci_re_d,
      P_W_rsci_q_d => CNN_main_simple_core_inst_P_W_rsci_q_d,
      P_B_rsci_radr_d => CNN_main_simple_core_inst_P_B_rsci_radr_d,
      P_B_rsci_re_d => P_B_rsci_re_d,
      P_B_rsci_q_d => CNN_main_simple_core_inst_P_B_rsci_q_d,
      memory_1_rsci_radr_d => CNN_main_simple_core_inst_memory_1_rsci_radr_d,
      memory_1_rsci_wadr_d => CNN_main_simple_core_inst_memory_1_rsci_wadr_d,
      memory_1_rsci_d_d => CNN_main_simple_core_inst_memory_1_rsci_d_d,
      memory_1_rsci_we_d => memory_1_rsci_we_d,
      memory_1_rsci_re_d => memory_1_rsci_re_d,
      memory_1_rsci_q_d => CNN_main_simple_core_inst_memory_1_rsci_q_d,
      memory_2_rsci_radr_d => CNN_main_simple_core_inst_memory_2_rsci_radr_d,
      memory_2_rsci_wadr_d => CNN_main_simple_core_inst_memory_2_rsci_wadr_d,
      memory_2_rsci_d_d => CNN_main_simple_core_inst_memory_2_rsci_d_d,
      memory_2_rsci_we_d => memory_2_rsci_we_d,
      memory_2_rsci_re_d => memory_2_rsci_re_d,
      memory_2_rsci_q_d => CNN_main_simple_core_inst_memory_2_rsci_q_d,
      image_rsci_re_d_pff => image_rsci_re_d_iff
    );
  index_rsc_dat <= CNN_main_simple_core_inst_index_rsc_dat;
  image_rsci_radr_d <= CNN_main_simple_core_inst_image_rsci_radr_d;
  CNN_main_simple_core_inst_image_rsci_q_d <= image_rsci_q_d;
  F_1_rsci_radr_d <= CNN_main_simple_core_inst_F_1_rsci_radr_d;
  CNN_main_simple_core_inst_F_1_rsci_q_d <= F_1_rsci_q_d;
  B_1_rsci_radr_d <= CNN_main_simple_core_inst_B_1_rsci_radr_d;
  CNN_main_simple_core_inst_B_1_rsci_q_d <= B_1_rsci_q_d;
  F_2_rsci_radr_d <= CNN_main_simple_core_inst_F_2_rsci_radr_d;
  CNN_main_simple_core_inst_F_2_rsci_q_d <= F_2_rsci_q_d;
  B_2_rsci_radr_d <= CNN_main_simple_core_inst_B_2_rsci_radr_d;
  CNN_main_simple_core_inst_B_2_rsci_q_d <= B_2_rsci_q_d;
  F_3_rsci_radr_d <= CNN_main_simple_core_inst_F_3_rsci_radr_d;
  CNN_main_simple_core_inst_F_3_rsci_q_d <= F_3_rsci_q_d;
  B_3_rsci_radr_d <= CNN_main_simple_core_inst_B_3_rsci_radr_d;
  CNN_main_simple_core_inst_B_3_rsci_q_d <= B_3_rsci_q_d;
  P_W_rsci_radr_d <= CNN_main_simple_core_inst_P_W_rsci_radr_d;
  CNN_main_simple_core_inst_P_W_rsci_q_d <= P_W_rsci_q_d;
  P_B_rsci_radr_d <= CNN_main_simple_core_inst_P_B_rsci_radr_d;
  CNN_main_simple_core_inst_P_B_rsci_q_d <= P_B_rsci_q_d;
  memory_1_rsci_radr_d <= CNN_main_simple_core_inst_memory_1_rsci_radr_d;
  memory_1_rsci_wadr_d <= CNN_main_simple_core_inst_memory_1_rsci_wadr_d;
  memory_1_rsci_d_d <= CNN_main_simple_core_inst_memory_1_rsci_d_d;
  CNN_main_simple_core_inst_memory_1_rsci_q_d <= memory_1_rsci_q_d;
  memory_2_rsci_radr_d <= CNN_main_simple_core_inst_memory_2_rsci_radr_d;
  memory_2_rsci_wadr_d <= CNN_main_simple_core_inst_memory_2_rsci_wadr_d;
  memory_2_rsci_d_d <= CNN_main_simple_core_inst_memory_2_rsci_d_d;
  CNN_main_simple_core_inst_memory_2_rsci_q_d <= memory_2_rsci_q_d;

END v18;



